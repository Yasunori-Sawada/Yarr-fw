`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
vVM59jSI2wl10h5DVzmSFIu7J9Tch7yqe5gFW1kFvQlrBZzGn6xOJ55PHFCgD5t2Bdocn3ZCfO3g
okY2HYdBFat+jfrF+9UewcJh7vOwOORXa3X4qSQvIMZvi01flNH6zm51Exv5Y3DLfq40ur/aFKiY
2D5QUDsNkNiXHCmKFEGgseMkjYvTQ960Qt3Nb5LLQzr/tRr4ueYMpKK8SAA01Q6iWIH591nfB8t7
g8BhDFQ7h3tm07/AGy8EC5MSPCFxRUnAKX1OYe1SBprX0ZKw4mPlE7/iyVGdEX9afwqZCAZ4thDO
K7BsXYtGVOG9UWjVRcl+AYR+0R8yb7ajndeJgg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
a2NZHEVZddQmbjNrJRh6DaFZplUtGtiVo953ZkGzGY/pQrPe5z9g77q0MjIfBzP26thVGRXsUpa9
N5ybmXKiqZPgq/RT+X1JsrTxp9/RtYc/11/sJnivazPjaFhsl5L1FgVLIqblqn/VzhX8DpZlDtIc
+Yz1ocoMI8ZnVblp9zU=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
aolUmSD8U+1mlCsZNX5xY5wniea86ZR3IaiFTGwVWq0Q9rbsG5KveIw13JQZtwvJbTHkyspRYe1W
yul5Oie5c9MO8PulP9tC3uFMd3Sz4efSxWXmap5FqaXSaDrTVPkmD86WAm5XZccoWG9QyXZkwEU6
YX7Wkk6YSTpyoX4Od9M=

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 250128)
`protect data_block
2jLmJV9j5HadfmTIcSC1hv5njhUC/K302U01BetpLv8koZdvpEKYHEX1fxACdiSbjkFY81cJOIs2
/dEKSD38Q0N29l7YCgXoEgpOvMW5SRKbvSf1mLtS2Cp9WVl1tMdqlP3fJtslVz/juj7N+UkvHZ9W
+toXoqMzxScPQttf7L3tA7Q6tcG+R82PiyYJwKT3nemmg2qzqbv7hjzaH5VPmqMhCwNd+Gwy56it
BFu4p6qpGK3TQSSNRzBvERUdo3kB0Sc1nGIG2q4K/Z1QSY0E6oIWy21FZ+LzB+tQVOsDU31jAC9w
/cHk2DxYnhruK+gkBN8cHXHkQTRDROIuGwgCg+kjv+/i8BAlfIUuG34N8Q9ZnsIZQXCxdq5AEdq1
nYIT7ovplG5WrVbkSZdqhTY7aSkgmnLR0OIUW7JVo7BYwq5Zy8GM1WP+HWCWmxvAiJTjDaHEPlqN
ghqo6alX0WjiNq0hONsx3kXOa3qKE6+A3//Lhvo73n1lSQTamnBHDL3eID66rHUfFI9jRnzSitps
ya53fIuLIYYtxjmHwEWdZIP0ZXb4ymsJEwYexiwkFz633lvJ4CPeWz9FrAtgvHi4U4OWFT26EtlH
qSLwZpNg219Xtk7+NdGKIJSZQW1EwXjzD9M4GooZ9xLKhzF+wcGc3lSvDVVXc9LBfQulH0conHM+
agVqbd0nRbCry7kmKkpngNqEhbC5xPFZmkMNg2q8jB262LHfIIlTzdd/BVy+4wT+aGxD+2vKu3lG
NAUbagpDGJ0Ik3XMUx+OqBQrd8E8bRSuBVkKGADJsK88F3k1YaSG25cGuzqAWa+tZt+Va/BErIUF
2dt4tZnQGoCj0+p95bq0gj2aH+jV7UQMDOsunSpGtqbIxIvpkEttxLx2Nd/XnNhYE4PCCZDbUny4
2mMiGdv7QkowBhrX76xaASdGhyQZM7/PGYpAuEozN0oRxatCY0pQ/A9G3ESpY8VtQ8+jk+uz0clG
2CV30sB1O+mF3acf9HVvwEHB5wIcLnA0Re2oWINvjqo4J34eLy3X4EONi9/SrgkDDn2H9rT9hrpq
CgbhD0tYzi2zOQFh/l1J6RFycGlmidrJ10NHnBSQ88t03WGbMJpBJURSYQMASbhJcgGNfPcoocTd
HLbppwhjqdp4BL7uDd34sDtGJO/YHkzvFbcYhwkB5FhmHV9yDHijxCiHyOjsBdZNhTD3o5qHsphX
9cf3E48PZt8LVAZblrz50LwhRMlzaQLzp5TDFEcM2lYTkx7ZSvQ7fa3aYFHCddXMK5zU1CrZAbmN
sIRhC7Fuo4a1UnPBP3zXFeMM67Cqb5eHunJCZW1ju+CB/Uun34Z+V7r/VLhsaKCon6jIV7tB4kvo
CQPLrRUpTO1INZQfXWhq1esoiiLaIxuVAMMMMNIoQRqUPgedhDZst7BvtW9+ApjneMZtpq9WoyUX
VnjlQaOeuOq+lrbX9bvhNUK07EuYxG7goQkynHYziWHipp0e8N9OKQLMYiYuIbrRQSLU0mwoOeCD
hskKjwGcczBvod6dcwau39Mawb4WZ7nGRZUH0o3JKMDfvazNzegXQAEyICNf/BTZJWj9jUXLvUMX
h1RUqDTWPID0i/drAJ8p5OQKQQwtEPoNNn6Lv0eqsUQ7GlM+jYWGQ/eZXw0ACNppxM56ZbuIky2q
OSO7o0BuarqGxI+5onuoBBly0pDKQO1x898vgEfXvrpZIw8JjxPKLkwV6WvJjytofPgwbtRMbB7n
4Su1q7b/4zzxNSs4gMgGlrwV3PYzaXmpErdDwBkiH19e4GiwP08EW40z9SduXTJwwHvRRocaigOv
9vLJJBIhrYIBqP3SYmiNnixFUm9uhS0hFVSdP7H9MKhoSmFr48Xs8EA91/INPW5j0yRvTOoMTQ3E
PDyOde3Ri5n4Khx1VGOm9O6jeYOLkT5RRxA480YjUeVj4p73gzTH6r/ByeRQHHU83Up03i4qN/dr
LQqJ2tQcA19mALqMb/u3aPvOXfaAftVBu0pO2JxX06QcEF2jbRPf0p0p/oxiH2wz7UlajmXkixMs
Te7EkjPWvUNN+VfC1oLf+CSJ8yDO/TXoc2uOAw6HBBf2DizZXg5jfu22QdyjypMFGLrGcB+rqDwz
iUlVGK0K4SzhQZmDsrB9zRj2sRp/v9cEqdRSXZ4mK2gmPgMtkO72xbuYTkvnn8OvaRwSRnDqIVja
BDvWA+57m6p1gJKySKIZNUXo/QWJVB/Vq3kfQfmWhSsuXuVvBP5K5o1TExxwjeMsY+R7GsUOyXFB
hTRYrB8pwvHmDFxbosU3R0NPugEDbWe16MV+j1X0o8W2ViexSWfLiWyy3vegBWxzItXRPEC35A7I
rrBcS7tfT8D6FFAF6yEawmEGrQgJtlUstSlOiyhkXSVVl/I06toKeKgktqxzCBABwnFfNnfkZ45F
ASV4jGjGQpm7rVwQRNE/UmOAjQ9h1Sa3k3WoeoLSQaYewbHT8qN9ZXP/0f7AkKmfr+7mRZYuID3u
vqDKGQlm618I54g/XDhHU/8Fox9Ln5ZisnwBzr89THCMRULX3n3G/PTfHSskvMsmkxeIugKSbeut
L43mp1YQsFpy+sUrUBO+x/BWDQmt4yVvUMXsu3aZWO/snAzDJfUiW60NHyEg/fKXV8+R/r28bVcd
LEqxm4DFUjyoKN0O7ericHdajt7AQ1y2a4Ocb7SirL0/lJuV9pZecdYE3cTDRr4EMnXCPdNu8rtB
dP6mAsQoZ3Jc8CAWFamGpxoxVS9s4zTgahD42woDc47RNhNsBhHAcx+ger/D8qPuunXXomy+mw8/
Fg78gmzlzcg+kXRhrxYdc4DBZYmnhlIkjQAZn6NGZSDj32JxNQHzZ4+xCphLdWQZK3oNWDgQmkmv
JZ6cq+pRsJIduqfgrOWnrWmlqzfWAxBzrx42KjYcV3ZXShiJv+cnUOrsPF45tie3kX20dpAY63Dp
uOPtnkkLNJEK5CraSMZO+pzv+6OY+gJlhzCVN/qqHU4V2DiD7QiHxR8+/q0Ctyb1ItzWcQ8FdCHI
d5DRE0S1k0sOh6zl6aKFNWebIEkn9/yZCcdlmFjkUMz4c2xum2B6FfdhZoZFF3zZWEJFpqUEyWdV
y6j1CZHIYfETgzW2lOZtQqmAMVFdL8LIbpiSmglyRvtvz/AYk7voTUl63OaIe9gcwsUHZk9mSZsG
u+jsP0ZfVXPmmOpXAFCoCFOpW1hAC4+6UBIUJKaIpiXed9I76TXsQpSJGZOFLUJcsKLVET3TY913
RuqOo3iXXkaenUnNvheg3f8wxNxox5FL9mDl8m29mLf+jO7LJQaxp5M/VdsjYmQpIovZIxD8pUcc
gnxkcOktaz7EFjAE81YDUkAkINcWJd/epqbiScDBPa8ANPbTc1OaYk4fqcuA/msEVHDOHCOzw8qn
8MfdcgOOJDzd81ebWjK8ZEuK57j6X9/FJOVIB8dp8vFSoyfbY7aOoK+/9ihz3hIppTUZtP5eqWzP
XXlEVjO8y3q0SlF3TIOgH5MGZ6skLh2vZSaR4u3yU23QP+U7uhpe9CdI7SRdG1KZhMj2lD/bfbLT
Opm4kWDItGq4GejLyRTOjF2ofl9+ioHh5Curd1Wh0ATPN0yKsIstodH92ppDjy6bgIR5D7c3WZ04
Zkeo8bXZZlDiZOvgoDE8G1kgm2uhokX/wQmqzUSvJQdMWpW3STOsQBZUM7vieLOpXYSDhdIuH3vy
omR3dfgf+4b2nyIOeiKLUZ4WabVlD0WPMnJzmJ7hwPopep7OZJgvnRy6Ci1/9PouW2dRyayLkLU/
FcK309B/96VwpTTpr9+U96c7x6n/jTdoC8FOONGRL6TPiuux+BmkGAHG4wOL2LNSOC2/4kpZPYCT
0Paw8pGkgwszzb7mYxl3npQn4l9xlrc39PnoczckQQZxU0HGM9uFqHNUQoofHG8bqbCuJDqPEEjp
sdiuVEQguv6nNhAwNA16ebLm8rAvhXHpw3iGF2yRKRS8dQK1hX2BTmgmtxG8wpyR/BCLt7k3mshV
tiJqSPT+zb3hjVl9KR7ecSmwNwK/5XJmRt0nQ/XB4/T5lzyOMf7CrKc75CJIWVOZem+Lz70r5+Oc
B4wP7I/FICdONOkvw/cjXWIM9xIKRFo6MfkpW2lVpe8pKpobSAjhIbZaNOWai5OEFLhfW4Ihh0ZD
wv8oGtYbc99qmofga9deSCnXW6YM69fkCTCApvxpNE8eqNtQoJ3NeIiEeVJR+0yT1q57QtBEyUh0
YCakEXXLUkOzWSTqiIpCsH02EOx/iMfYGa8ck7IkzdHrVDjrh0ySZ2htXl0Mnc26SPHRW7cD/+WM
u51l38g3s3qvW1VnitEsIz7SIjwjbUZNaXVF4FpG+D5mOO2G/V/RDTYXH2WIdDUM1uVZ1McIIsa1
CoUgiy4q9UQdpk/AbbvW3VMB0RpblcTLXMpSmwJHCLawInr+qBgpnMMW7F2ffdCnz3X9tZvHcfEu
7GgJFC8xWnOuRXZiH2knK9KnK6AO3rrSKaYmbYZvmIqvA0AaQOItM8wGiOPKWik8xuSdFIobQuoV
U/eBagoiyBMi/hVTKP+1Fm0j4AaIsuzL2WswuYp4+9CJIJf1Av55vZNCUQZpSvvADNt0bxEeTLZo
kseW9O/BZLaqF/KWZ+LpFdadYZwUS8pDiqFcbgZYA1lTlH1w7Q4zpduUVzqoCz9LZScnBI052+YZ
K5gMDSER69h5y74SJ2rRalNveTTsDYlvy9lOaU/QKWfCTX28/eGIRrDaAzYwXkfgxHm/70CLY1Rb
ki6V7Pg7ugTjEFebsl2+BRhwiCpKWR2NVAcbBXlubKQqPgrU+8ZNE/kVcDIwAzESkk84R+jUqOhI
XU8930rjs3X7dSl91NWp7FFxG5jzBp25BZKZcAym/kRsjuDyAD8wjpCT5tONp0j7n07BUiRzY3qf
+IeywWAIesBNxwDxZH2VXevHMQs2dbPuz2WKXGg2NbXZvta2n09se/3uZyMUL6569k9J9c0Q6YWx
R3W6uDbTzaDtWo39CJr8xmc5B3nNDEeWMD1gInZk7ZA2WgOU8KpBVQZWhKSs0lH8X0RU1klqp2im
XeFUCXOnij5ZPTdhwYCfLKySBt3zkDSZQa7K5zmZrM3DjNeKRi7vk4gpN1dm1cQpSmyNV8mBQ4Mt
XM8s3gmEuIoRYGY1CUpchoxjXtF0gMx8oUwpmQlO31A4q8vu1a+SAT3Ibo+5vy/EU6ekJSXAJ2K2
C9wCOeO0hW0hKEedGfOez291H8vJberAuKor4InVF0XlHglsXJlGdpRgjXft/7oBkhqfnf1ykbpo
zgXKfCBWbMOamb0qq3h0m3rrGA4OQfG54dt2KIETcn9NxmOBW5cvpzONXT2o0SvN2M/jr2Y5jcYy
qmPC/AYD4wiBZUlrnYw/FAZ6o6yJvWGITjlrE0Wph301SyZU5n1HeOrVU+6yGDKy55+OtuQ7Pjd9
KGrKH0MBZ/9A8fCMA/cRBHYmNfNprexwVhCgC4neFIg0X+1YZcy0FCLoakqSi/ev2QXy84o2RdFo
vs7rrBo9JSJ0YGRnNMfJLMlLEZx1uIFmIdSDPeHz6MI7krE6eCs2zxZvFFrlx5flIiD0hht8oDpn
UKPCBiVA4wlz9I7Zh1YShrfb2LpbQib38FUc/gmRgMRB0P+FPy1lIP70p1ZRWkdBRB2v49/5+X8J
ooIgv+FJ6P05lZofwD9ickyVxLOTZCb4Nd+I8tER2J/Veo+bD1JD7CzsArdp035myfdrAwg0GBOc
6eiaV4DAmXT2kDMb08uHWQL+BL7vwD4D+hBsapdsATwCNr1V3oG4YlHOjW5eC4tge7N4V/6VPQmP
WA6mjm/pt4Kt6Mn3rv+Q6dIzt2OdLsCQoIigWp2p6Ey/x54mZlPHR/M0baFXrWSk83/vO1YmHdub
+hoci0eHC1+TMCDdEVCd85swNimPMM+GP9yYyu3KjsiNddKzuc2GAUgWwOOA63dfqPlvaRH2muVe
QT59mgeuvfcnyNJqrnOuzMuX4WyUChKZxp2YvSPFQRYvzzm2sbjXrkSBplJB8ED6VGNEb9QaugWL
mc1FivEmlE0K0VWiG1FqKQtt+dsY432szO967zMAoAhoxWYQK1GQy2anf2XWRiC8WhB0TZQtoDJX
9nK0lorKGD2mZWX7egwKP4x9/LFAg36qKpvZyA7XlKholM2Lv/dE1tiUfIkHnaMId8DmhyKRhUkj
ch/wX6vcVF7coQJxELwmJe1ZWY1N2LlGm3dny2j5t0sD20GG6GE4tjM9jka7FA5JRGe9oA7ZEYy8
+bNsqigev+IP/ONvpjNsJXWBNm3PWQfK1qS6eyg2Ct1by35bWuv5skr0vxf3QDoKkgn2f6rB4hdy
9EXHOIdKDA6dRw17cxN0J7ilnS4w81yEL2jqrfzM8zwwKy82JbWZ152TS+41U8GasSsSg6vU/Uxr
p8/PRn5jylhJ/XSOfjbbgDLtqz+0S5N3o5QCaoIHS5Os15JGN3FsQGzH5ai93PNFg2rz/IXoHIEH
vRqEATcxnODlxNDyKaA+AA8HrvN/grMnVA+e+awphm/cZ8U7D8O1dB/WkuJWAJJXb8XVjUibDtuY
EFQ2he28nR8cxew9NW7G7bUPDYO0YDmgc0NjJf2ew+xmmEKFSUXs80i4ygFL0Ei/x7bc49TgTn/F
EZY0nhSM72PbMpdISUZ/IXE+/uzW87ZnoFC0dVO2QONWJYv2TvCHz1QIXepJZ4uc6HmS3ocPrYNz
xEXjjsYCPa+8MGG6v8QJrBKlzeaXSjiaMBAMediwHWrAPsp6MYgV1PrktXxS1tyO8lGmKB4bgqgi
6TiLHd/ju/L67j/tUTzT5I9WQT7r6cBNbUuSLRJI/UQ/pDg6Qn45Zr2kvekhF258quU9e+GPyvjR
uezkzFZxAlJm8v8j44carQBX/6Ea6xGFFPCHWvVQPgv4TY6Y46OXeozHz+cXKevkeJFsnGDyUbY3
o/8DEsAjoq7/yjDIZUyQ+t85WrbtP4Q5Lk5dYYlHgsgkWyhayq2cr67EtEwdEXGaRS0Hn1OAM367
ZEAc4S8BCD8wdKZd9EUdrpCucTyXvO9au2qcBNZIFQM4RNsgpUeDFzkB96PQZZtL8p0NpWTUnm+S
p/TToDHHwzhd0UTa647c8Wcz4aVFxicPxVEgDmBf7yAxlBlhQLdw93HwxxHjWB5QFF2L16phG6Lx
gq8yVkCh9Tpx/+70bTcFH0hbjdknjeCge2z1qmzKuMdCME0CXTBpHwFjy4PCD9LLMw9OamBkeC8d
CDRwRJjqBvxAenkhcXy/0uTYoqEEdLh+DHTD8yP84KCOAVcKgvdaGl3yQyBvKFLnHHoYAVZFFAWb
/bPhXdACrcY5mRDuIwYsitv0q7AFHoklZfYCENQppX7rhi4ZtEhVLPoKGAuCTwyE4CpDRTCo25j/
BfTrbipDAcGiRKjkzXEJNnTTaETHY24skPhPfGja/2C9PvRTrESrsdnwHEHpweWi3vyIHH7KPtX0
3T/9aA+LveFy4CEy7yAeTHxjnCtRc3KqeKCdFyukLX3pKbnXrWr18nFufEwAAS3k5HeoDD0/puSV
4fM5yJ3/cCB8wwoMq8Fc5A2cvDRkd6LNjGVMPFkFhmeXYXeQuAtfPer06SuqwqMO706kislnl1nb
vR9Yo7Q8hpx4Vnfepb/uw5ppPelcyDOiFbcqCJO3ccuyEbBeEA9lCRvKsIGROYIeCL73FFnjAXr0
5+iLZqNTq3uE4is5gNXdhy+pe8zdBYxnubPGQc9jci/S9pPwC0NJpRNX07a1zXfxSNZq13QI8hMb
qsAgNpwZZnD4Qb/WYEA902viLHS6cz7IT3FljS7UhrCA0/kbjp70T04D0TJMbkG2ILCqZ9u50s+C
eGwoKsI2EZdeKdTP/iOoLZ23hIo4HFNm8oC+4aQAXePkYnzrc2OsUOVU+X9TuE9SldZhx/McY9hw
XDkSD5QwXPVRbjEBvK14qFNX1LmjesKbvR+lfzfWMRURx5WfOPtJQ7x4qfW+AIHedMxjxUMNPYk6
8Blzg5dXzl2EQQakHqQLKTEsLrNuWN3HFJHdu/OEqAqsAZ/KKlfqBTTik4XFnNFJ4EDvTdSA2swT
XtA9vdrZzo/F7T5lgbdkuMRnX/ZmmhICifGmdzr8kbX+u6IWtEG7X1zXXglY4X9Q/0zajYePnAGk
xMM8Asa4ZOJ3OjGdmuTQZFwEozYZDUovVUAcy7U4zosq/pjzYwNQqr1XJE/pjbo0hqBsXGqSUWJM
iFbC1yHkK8rQmU1AQSs15NALHy2eG+gdEuBkoTTbtC+nrnls+NCBAT5N7k3EG8+B57aG9P5Vsg3a
MDljrvaa1Aya+Sa9egtuaotHn4eVT3xZLnt+ooxXVIZf2LAZrzA+WqpGxtWM4GV53sz5+r117DLI
m+yye2O2btIaEvmPVe3QiKFSRF49ynA0jYexJzaHQtXCotFCoJNJTWDV2qhz0tCWq/k4ooW6Kkgw
r9rQ/kKcwumbDEWWcA6iIeVJHasmGdAt4No61Aw0B34FNYcbU8oFHDlW5kM0ujkH0YxsWOlvA/9j
Y+lo1sZUfH53i2jUi7oXe6Fcup5lz3H3rIF65I+bz6CWvscza7p+XePhZ2aek1wzJGy1TEu651OJ
NVcykwAOAS0cZN8EDZwCl7on8ebiP9oJachq1NjNBR/XojX+JWbmQLxKbyMjo94Zi3LIEVTBSvkZ
skp4eOWY+tGH6nGPqwalmMtOcry++5UrC1vxB1K0fH4N7/tkE/lpma9hKOa3hEIwB4PgoxWoClIq
XhX3/7XqIhpL0g+eBHBTS7c5zloK+cz2gUiFIRqhxCSkP9i5D7fYSgyCELLDKTFzIh1Cunl6jTek
z/FW/kxQ+EcjdZl+nUoN0zY5DtZtcvntM4DqxLH1k2/yU57fNSxHVmXuObILE3crjx47PVPJ88km
cwJmPizRym3upabZzjFG2W/RC35yZVp9a/c3UlVXdHsBMSD/DAdPhFqP+81VM2RW+uiDXTqxLTDe
aPIcK70cSowEuDz9cGeCZLWb/w5J0ZYoEhnPKZPF2RZRg+eU19exty/BxD86c9EU16DsnkF1dEfH
2M1CK7CgvXgrTVLIG+M6MOgS8J6wEYHd14d0dfsaJWdGQh8mmILNnPlLS0ZTnpdI48e07RAGojMi
RTrjYw4mLcyzGS1wgCnHbRBjwtdD74Ok5NA2WsQ4+Ebqz8DS1H7wuWx7LbCW3E1yzg1v4IYU5cpX
mbnNaH99XUyYguQ0B6kBgWSi/+ROFtjGwTgbgbvD15mwFvz2t9xar8zggJ1wsG4+Mo/XOmOuuEU/
27Ic905LePXlKnFi7UmYTLtaOA1+5MotueDyts3S9++pFKt7MuEOwZYv5tnsbffiSW8Y5RbSY7fC
XaNqTKEvguGVnz4q7xBU+nMbzJle6EOQOgm9Qr6cdoevzDg79w35HyYMN2FsmqoqHvXmr/MdODt6
wmaCzG47G89VUq5j+UjZqdv5XuJZYS3pcLpMYCiwT5BGk6dflaeXkfB7q5+zooKy/4eoGIMfgQeg
uvEXmzxbnK/g0M2JcpuWuxYpaWjsIqXYEPfqZm1rasWfitwpEYxldIrWOMmKSE1hxmVEjgsPjT2Y
je+3MQZWiY410e5ctffNcHANdw02OdIszRSGqi00Ltk4b8LNBakfPHgdsXILBKVRv+flcuLcBsaS
yEHha03eEDf+hYzKh8JcK2gdB4AWbES6XGKHHLyN0YANRGOs0HV6N3G3e2FP3HI67Gv71X+s7PA3
Ui/oXGtJgmdO72Ey5AYEtwh0An95m3NWp78+ws76kihq8LFB+smbT6QCrsHjmcZJE7LzSAOd4Z2T
M11L36G2c7rDEZX+cS7Qi8m6qroGD743Q2LDPHPwNQPJd9GGt3ypb97uV4ZuBXYyavbZNhTLWu7p
QnO4UdEpkWPiKP0Urc8tta5UwRFCH/5iApGdlq9vItkrG7xjfEDOp9G+z8vKxfcZgqXlLDAy071i
XxYjHRNjXR3isEjGS7zA+PEWdfYhjJJPE9XZ3778TUljcIXHDTUPd0WCiX3zU7p5I1bgwWp5iOfo
drLiP6kEGtVyyoSFoJSdI0tlIM3UxIezUayY2+zCvhPyWXnp4OP8PvGKwims7yVwffvbkuJpUu7c
NrKWhWikid3PlHYmqTn+l9pEfiIy4FIYqrmGAbiB/vxamNwau0d/RDSsB0jrcpajUfqsqG/ljnjX
qQ6BVqRp3MIyXWT+rn2ws5X6JvfzWKn7ozwnaolyVwCJwTrJCQCXwd5rNclJPkZl7mhdbxK7XZVD
QZvB20UfarnxCOmCFV1JmPuENDq/Jwo+NQY1X1deHnvzmjtHdtremmy0mLDBj2rD/hJj/OXAKuCe
ojsOxjRVm3OcMDq/K1J2tjVhXcD5h1gn6k5F74qxoJvYN0X1t1ZTY/suni/Jm6QCGxKMgQt77/0G
FYMTn1dEhWI6aKD+QfJHwX2BPJEGYrZFVTRtL5LIa8zr1oYSUTDt7e9eorsqPxhfMI3JSIU/706r
hK7yDXfjj9MxKwvldkSwyGaP3NvcuT8HHcIndLKrgG8DXdXJczrp4VjrZlTTWnI+F86pCxdp50Sr
E30Tyu8q/OAhfhIF9rtXW3IrFt47qrXEfLaCqAe1vpmyxYvDMpNarcS1Ng0lMoWo7BNym3xJ9gOK
oXuuZ1ZHl0unBEaSCuCEDiP1nUXRtlvmZMBa7J7tBLrNyiz4+F5bskx/CT/92Usr+C94IHHBJVSH
kjP0+AQY4Ng+BcHH6+HykPcDjSuDkcnsOUcQ7PM+Xq6ahL22TUOqrIZE1cLbOal4l4BqO3sG83RZ
E2HrctH9IbzKj0bTmRwCffskkaIQYnNMFRLtJw+oU39Hs0OaiHNHF4yRhZ6rv3FGRK8OnfsIJfzI
FovlQ+VjBEFBJ4WNz5KwiP+lcnhE82xXRwIX/UAwzkMKPev1T5IseOvDJ4253ZJs2h59wNhiXqK0
2CVws7AKYG7dZ0aPB70LdggO2bhlnlzNdsQmcvZEQgH+ouoiCr3Kl0C80af9K516UNi9kDNHONLh
/vBZpKWEr3accUKgxGt7xt/bnZWJddQ1SmHQubN6HPiN/nz/OnMVIx6Lh4DIJbUQhp5maqOSaW/D
qr8p8gNOtD6TW2OGl2b98F1/HZbjgBnaRpiLABk7dVzN6sBG7bqn5/4JlH78FbSpMLrEIosDcCNt
CQMqZdWUT729VNOk/J7qGP//rPIzFsFWHtsGTJPOy9Lz4yOEGbR/3oH4qsxqfsF28vF1dkzIShu8
4E2J9FB9Ib9JTuVUHR8b6+XAQq7s7MTGfW07cXe+O3o3h4RY68dswELyYwQDKz+KtERyhbQ5H25L
56DaTwZMgXXyEAGIIrbU+MdOpZkMLSxTZc1JGd3mEnWGW+M8Jux128Q5Ru/llHBtt+hnkzA3uf5Y
lmrRNfMKfL2qJWNOyQhDU0XRA0P12+M1K6xxlZ5tpyuSK5nWKcoWfmzWuZI6Kb4jb2wwGk9vgEE4
CDg5kNAH2QbaBAYGHSnCTjXnofRkkYEBXbWAYkOD8ZclM66rQilXNuPlJLiOzQogaj5wrLeMQnvh
q/+RVQJnXpPmCoQeGM8+aG68wT3uNt9gwj71IzjIYPCi/tgh4fr3b3WK1Oj5V/gJjCPIMhVg5yzA
GT2U/rANuLuYQJO4kskaH6mI/zWQV/blKcQbVh9akRaUoTXzgvNVzj1U53kwVm7DDG+grpG7xQBs
GYQohG+JH0f/SR8M3+TS61c8DpEc9QrKOCbHYPNPoQaLxJHFKde78u57InTOyZmg0iwAOEj0X+Zg
fmlSy2sruFIsF43Z7r6XqhevLppLmKAMzqYNggmDOE/lIaBTfdrqHEdl/xoNViZ47tsYWdcxyw+X
iz3q7vHJQIHb9YQUY9XwD2qjLGb4Ygefrdl1QOvz7UKxDa/p2NYLKajpl3SOZQirM0+grDzitAYP
UjrDS4R9QAezF/fyDrmcCKtta9RT9e0ZBsXTDiBI1ZWv7tKb8LJAZi7SxSNdCU2qS0vlX27WiCzu
iBdEHzY+6hbXZEJKPifTK5LfF+JnqhdRI+QKZQc0QC3WzXjJefj3L2w7wpvAMn+CT7S1vnemZCRF
eGBH1Tx6FBDiF+dj/44HG8WXVsOAVusJGrtAehmuV3nAfYlyl6JW8nT5ET4HQ1BnufcAC+Aspiky
LARDjASz2CTBsU4ZscGE2Ji0c+p1t6Q4UWPQv22jKfCa44ovHYm8AxqgqVZPLPowgE2z7cR3Y2bf
Zwtos0222oStl2UdRYj2CjNRu5AUAd02aiZ+BtcgoJSWQLCAg0Rbf9oxfTDqCP0t+3Utul1b4HIx
Aq5NjxL/hAcIH8L4XKfR4i2ffvN5zXjz4BFG5DBDO5q0/gcyiIoiVpnRyWMYdluWeCRkzEJemDeW
6jcUM4Ii2NBcCoB79F7MsU+MYd52nzj/Ve/r/bh5KMxSWR7idYqn0WcbMgjS0XwnZg6RhBgH2ACQ
qCCLqMdDiGy/v5pyd68kEfI1137B3zaygYD4BvYCqYYvA/ka1remLAeLkkn7ATMTEJC49hnZFXW5
tN5SARGyGkZ6he5jEdJ7KbPeysKx+nlrrn0+X0F6DfI22yzLjOvX9JT07IycNnhB+meWYbFd3oQr
V9Wpza9eZqORaSuK8DuQB90V1mFEQhe19ChwdlDRWriX3BnBSpZC0CGYhdct7y6zNNgMfQiNHFPo
PHN3Dmtp+07XtyTFMtMkVDx3pdcVHuMTj65ELm7fVU4rZZNm9alAI7/PBxic+3XNMtfvvlFoNFOI
BFSK+EcWXEd/46cNz7SflhUQrow5+6QX5K77SP9MlxugK0Z8xCSWnNtgjRtRYKXwlTvzvUG9BWC1
ET2UB0AflyLqcvMgvxDKwWmAtRdALGzDSwtBm0AKjhjyPJj0vhrlIay1OIzrk8EzhiawwV1zK8BF
JJ6lFEJUtV00yNMNjW1ewmHIYkaXcFmDH4LnlB+ldsvN2gmTiDbOgorFwi8pUD8ykZoY5uVR3MDW
45xIEZ0ohg3LaUvXViHk+1TnirgGG9Hnoq1IM4ZLmFLO3l8J39YVJLyDEsp+kKsCIQJoCmI/9+np
NAhYucM+X4jm+TEAew7ApcwRFBDmC8qA7xUkwE3l/hgRYT4kOshcQ5gb329p9t04a/T/GVAtM/29
lFEsJYxVTw2s5v+XmJy+qQNEEFKUdFzAbyDjCTRsA/2obrQrgO6JtPDM/e9sn2T0AE0uVN/yuHpb
ZEdp2UTwC1jqsQzfhDfZ6Wi4I9VEIqbPVd0uPCiet2SDpT9X68aRCfq3JbwtO3AcP2KAygPooxxJ
7qJ/Y+xN/C4AgP3mofgMX3rz1o+hilSgSXiT9o/Ht0dm1t4gJHROODLsmP93WClYBXiPEWfjUY7L
k0u1rI2tmGF3eW0ZJlOZ+m0VkRf3Bplq4qof3pMnoOQYK0g1gbzvazvAP+8SG6cKTykxgInsDAin
CkcEaxghwzKkZ80ZBr0EDZYbC6xWHffvIJYksEktJ+RI5Iw9rR7nCmpZJGpyIw0zTFr38d4ta0r5
ZWhK+3XsQARKpUAazkv8KE/IofUT3PCZyLFnFa4icYhiAhoYrZCY2XvvUNwQWD1WEjNr3vhGrw6o
QU4cMRISXSkBXSby3jOozCr2HcJRkpD6cKrvxscy6+imqlf/xj0K2qCbGlNmMxfaZFtO1va2f1A2
tfkm566TNrGxU+P2ZlDx9A/d0P3i6jEH2fCgVTCLlAn3dVWUH1d4dKWj8eEiE3hmvRL5UmYInznU
9C0BQ6WpKqkfXtcN7eP9OzyllEAi7h5f52PYnvRyYTlA232zT80lhZMhgV8Qh9hRmJ0aT7bZ1Oe/
pQagPawKP6njV/jMNmTTYYAxidqk2X+9hN2juVZCdBXVWu471OwycvsRUXbjpnvdcPxv7vo85cDZ
O6q2KsboVYaeTB+6yelo6IlI16pTNxDQ2bF2LzG93i62qlhunVdcRrJfSbOYoFW+BJXorZ7zyIco
2N6BznEMitK/G0MrPZsyPwXO4q1Me0w7dWzFdoqiOu1bP0Av2dkvakPA9R/PhN9aFOZO20PCzEvR
WPqCzXOA4ew7inTz2xb+GTulHNE5yqM/iWHNaSyX0SAXlDuT3XFjpCPIk9n3SoWeWdxdwdo/YSKa
KzRGR6owJuTkKk9ZOR4Rs4chG8bcUKWp5toAHvDdXjCRkCUtvsyUuJ6y/Ik14sJFhb/3KywfKoxk
Ye6spvqcKV6hENEnpyKGlT1kJ+yVoIOkJJDqT+yk5WAxzTBG+EfWmLg06x/Ks+FksZ4Kq00X48nA
FbS4bWKF+ajOE4WAvWDweJk78t0IZNQt7+knWd0L/abdXtbVc0619dnEUi7Ji+LtjDIRdyS1rJpZ
pqfDO0O8EuxOp8bR8tY4S9gIM2N7b03vEc+O0BYPZhloWgEujdoWbD5JWByu8Kk/dJFhZwgzIWTN
661Pdn3THQywHlZI6THz0Q/0ulbYPANMJ4ADj2KRctwQ9wgElejA+Y6idmiVgCZ37odPnyvjLAfn
DWBlhlSW1s8DOYXDh5vhAA4jvonHU9BBTTfeZRI1qyCIXViEKebUMjozkuF5S31ldfVR0WyT3p2o
VLSj6GFz3vtEUMLQvikxvjQ0r6dXOu13Y9uMYT2VjVS+4AxM+7qmA1ArFoApqAPUNEdkJJEej6CW
ipxAd0Z0CiLa54Oj1vRUI9cjudYNQPZH4qSuiRy2/0FVKcO0Y34HBDjqPMTXsYtCJffrisomGpUn
NRFDCrAydAv9E7Tiec27BFDtloXceQksFc1y5gHpO1m5j8yAO+QLdE4G1Kyi0IbPTGO2BlaCGg2I
lraKj6bMsbOaGzZi6rhi8btzZLoSThZ5pfs3vmYgVFD16d1ISHqnubd5u8E4603pQAeaecuiCS6M
YT9KQAUM8BbJ9xdpXI9RwUDKsF7H3R+fhwClWY/KEWrcVnAOtIoGi0NianPAmKY7F3SG4yr4aARE
aWaWN1s1RScCirEcrrjzUeRY8VoM9jH/e+n5I1vu/EAJMCs4EfQsLQXSkmupZ+CTuKuBlJ/SF539
0avS5KtnFZiqURGB8BdZNcnDe4mQveDBf25uxHjylAj4HwxMR3SNU7JgwLo46y5kLBT3menLebEi
xYxBwyxF9872Qy9R54u3x6wj+54+/y8HQ0y2MA6sJw5GZjMIBeZl+zigh3r04bgXHVCXX1sNCDCc
CZaWqojzlL2TMNBn2jbLJg4ueixHf6yZiw4kmj7lHJCgIx3yW9/P6em6pBSbvQb+BVx+Ujv2qKXk
fQT3nIEd8d76Gyd0xHhTnN6WuUnklJhqz7Y6VIiro/pADa/l1LT7FjySUbriA/djOu9NIVrGfl86
BUJ1s+9vvoH2VLfkGF8daECK1cfZno+A4qNdcvgRgagv9xkUsHO1rCyL28ewU2gFtC59QLaLMi/0
lFWO4WN5iJxEc8N7RPvE4+NM7Zy2xALJVjc0CVpezi3sDcZC8Bwq7lVPuCh+miJIDn0tvQ9CEfkK
RZI5rBlw6VAItiekTUS+6qIB13pWrtXppgsBC2QqCP08Ckzs4p7BljeNWi5d8sQCfvEJPG/IQhNn
vFIW1f7R4jsdXIYzOQCYCX/kVftA8mZk/T11KoNJHSAxhRybxSuhBKWUqyILoWMJ5I8YfaTYjOl/
+ajtRnWy1kkR0r+seHXepN2cmifaB5vWqpycciXRwPQafEEd0xeGSekxIZ6VwZQPV9tQsG078BaO
KEduY2NGHcbSsDN+aUr3lOXJzvWtg8CiivWAbuIco7dM4ruKhBpspd/OozHkwSUgy/J/AHaCj747
udMIR47gYB0Kng8CNj715pZbwTDrgsgu2golfmx6uxdCG/D5YGowJz5csFciGJ1oYZPCkonySwPG
NVHiYfHbjwQzrYK++fe42jSx/QZG7M2SXZlTpwYUIw8ihSdkNlQ+XoAn6tRippr/JLqLjyEinRXH
ZBqj/5VD0qla1o/lh/PsToKIDtMtPyyI878KTP+1eteb+HW/aRvwo1fGHOtez910S5uRRNypbcpX
jhk3cbI1axPaDNXGP6TiIS9uJx/3/c+MglLBg0wOoSlUe6dLnhcJnAqWJh5gOw3Fom0/77Nt8on9
TRLr6IF1PKPcnh82AjodSaYiYwhGU0iqWROlYn4Oy/w0CHQJKt/97EP3mg/e3xZj5Jz6LRmgBueF
8YI9iyVxD7xuJABy5dpzRUSLFZnHOZDoM5rsjpT9xgzReXZg8eldmAIMalG0HpMPBs6ZY9kV9830
ZO1ky4ns+KHctlPMsW6AvRHpJZ525XnNjTO9qAOYzfy2VG6pA8hVE++SssY03CZMCOaRr/XLDoEV
/ZoBl5QbtFgnFTk0RphuLWjjOsPsVwao2/6/sRu6FjwnS6NLjtblcUNsqW7zTwYoV9imweTFRnu1
0sS5t9K0mtYZU61opwaUiNAeaQb+2YT0eIG5CqefpOP+aORPNQasMN7nN89dzmVemnzLt4pnosPu
IGNIVQ5v/Fe4wCjuYoi9S64RwreIcQxCt/0Mtb2UMnRBlc7NZgdXujFALekKVapvFw29vr4VW/YN
DNZtn5FhqRVjwye4NM3vsfPt6nHuhw9qbcMnBuXWFadY1fHFwjmONfBFt4LYDnZbbWrouCvMj2UA
/MBpVBXhk/d4c8i3z3vkB3zM9+5O4zsXyEOTro0qva2ZVaidYXdB6DOPOwjREp/owqQjCOz1fxK+
8dMCODtQQds5Z8kg7Rw/ca3HrWe8A7QBsxNXx6W2HFX9llW9k8uE54VWbj9UPeRNc1lhnvB6eUnD
E9Gdex+tUG8Nhp51IE282JFnSO/fLHzEPiWpMjHsi1CQV7whAnvqzBCCC6V/2aSN2jBYw0GAZIKk
zhKhYQc35tBn4rOVZ9xlVcmCyMmKe1Hfcu2nkimrKC919QSsihvzpz+8YmORUFriStaMdX/6vd3C
fPUojy+WG62OeW+whNgTy0acSqhrrqEESf4+Jre8gqEssrpMmObGJkpT/vDsW+s+YYN6lcj/ELyA
jiF973Z5AE1aCMgSHokt9Adtkf0BA79ccygHFzpaXwFyva0uYc4m2bNpVPI+eeePZqr18ctx2Jx+
cvZredqK9CDVEXByOOQ726kZCzGD7yNWIwfcbIjkJu41/5ENFkD8OFQha4iA7UFq0P/PPp5VSCIe
XUWUgfiiY5vl8TGWJvJlj/615aGZMyo6ULYo4QHGcChMcD1jJFS9mJZk7HuG6OgZfoSSLC0TXq5D
lBAUX9RO5aEeM7/rsqht20VAafdiJFsbqNu6KdEyLm8fMTZAUNTYaJ0sz9vqknye52jvXNYJXwXA
841EXBL82ze3vA6jbB+v/ogwaQB2JVVGX355rQ3rwyEVXME4QJVgU/5YGpjJBaHdSpBtkix7rtIN
w783Ywr+xQ5WtEf0JSYxean4fEXuXOIS/FaVWRqm6G1Y3XyupRbSKSKardS6tKGStvy6aPdVlcNm
McXJzLj+985oi59l0VifTt6sujt+M6MKI/zttYfQloDRRFpe0Ye8hCQpqyJtTYk4n8dkMFmrJDmM
wYwFmj+WZfA5RANMxFD1SsBrcmwRSQXT9bESZppaW4gTy792XnHyKOVKQJgfwLP3VWJqsl+US0EY
hOSVE24OsN5ckcwG1eEuDaynwgnqVQ1LJOfQNmyJuxQMlYPf8TFhkrA6yeIt/n24Mv0bRFjFPDph
8g2qEu7VDOrSlRO8aiPvncLXOUXBqHim6WyXv8Ponr3APRvvHB8jwb+IFzunngWkR6U9U3gTLk0k
w5vHfcv0g3bZfpRKuk/BEwdZxD3TATMSMonQGIQ4O5QIkffxVuBUsq2o1itSEY1x6WgPAN7eWMAb
FWg1OTCnS8Zr7DKrkfwtzw4npK9vbRRewuenDOLOZ3BEGVa7r1JBfDb80us1WxByVTgyOYOytWkp
2ifmwIlbsq+ePWoCP0QW1VupWuQPRQW88IQfpVY1n4xUgcbQwE2gBEg7wSRJD4u0uQYe5GprqVaG
eL7acYjZ3xV3T7GNW5q8N7Ecq6G7iaSujaXKR7Q9cSpBD4hMOJQjd53mC3XTtTfJrlyRI0K6XkOq
dXG5537jCLn61gWEnR/7TM32BNYsYpfnzqhliu2TowT5CQlE0mLe9VetwgPaIdeSErsM4vLKukM5
uvJ4+tiNYjemNVG/82uAGC2gmbXouGng+Z7MzA/pEs6KinydL+Qnh7yeHbLT5mHGBOGR4AM0yPEc
xxuHh0sgcf2EiqSQTXRncyXqlvcDjdua7FHFW4h5Fgzvw4PUABPA7pEUNO+BbWX83QZsyh34kTLV
hppWCDPmlU+BkTyPX5+QiGfCHbsKazHw2WnNDkC4EP8I7/Oyo8qkx17UfmaSrjRFVDIIwILKDcDC
UZxst6waCopEbPY1/AOsX2ewL5v/va+3EFfQiYqkS0A17E5S21q9rbcCiuogwOGz0AT+BkQ45DwX
hdEe7MbiaGlfAvfljb1JVNMVRBeulBsajAGyr8ocyhMdoXYiw7U1mAfluFM8JJliWsWtD2ptDEt7
gDdErWxQPEj0RFyXsXNITQEQrtnRvN9rWxlLxEBBgJtjNFc4BtaVuWiYdLbkvfCNSKNTPNYIXokQ
89Nlr+yOJxvWbTleUP90AWIsBRISIpOu2qPuxZnjQdqcWMGnZNoUFYV0TjGe8GLDdjiy3aNd8F/S
LO0oKN0fZdj5TD5bdhBOnI1yDs/lRtYE1LPjXL4skPBRgZE6KqEUOW2FQntUwwE13hjTVGEdVTwN
BNUn1LS6zh1x8DEUpXPOFnMQjHggLe5GmgHq8GtPpVqCkiBI5WjoERvpFCBiifBi0T4OaBKp9+J8
XcV7H0pm04+3LY+2sPQNW9DTaflhZWvSknAM17TTVBUdKaIASzn1r51tJPEnmG7Rh8XDsxLgbSXu
MeQk0OcJWs93vlOYyvvcj23FwS/Vx94fCSr0Qxm6w7/4VZehJb9/i+2gQKbzhzXjXH9QNN40iSIZ
If4sDrvofN99S9MThN08JpOXYU9Qys71CLQcFiIL0k+fc+BRtPMMWuaXvBXM20xhmp60d2xCYFgD
HSJWMW8GLF6uMn9Dvbzpv83BICjL7bcEaKfC13X6SjZFhnwaAngmpUqyBicZNMmXWmthPFacuYLQ
GROeQ3uyID5We4YPDlB5VXxnZ1QThCmViNj8RZLmDNuaAedAs3hDwEmlyalvZuPfczaXeqFZPlWf
QoGjslhIoKBQyTQOaihh10B6UIhfSbzoGQ4D6CYUGjELlvOpq/vPPT6N9sB7MKNsUyVt5Y/mG21I
YrlQYqclrV1AalFCMFWObCHvRJGVd6BqIjkfsM/AbBUsphhfypEBA3ssEB7WGcG/VPe9GLjF5crm
uJBJi4PYo4KXWo+hK6N2Fl499BhKU2hMUt/jUPuXquAOf6eaJjGOp1bbSQ16L3ZsmbJnA/4vb7X5
Ad5KF5RlF6Z41S3rxwWlXrBAouz5LOeO6aTPkZNCj69bEM06x1YdmcLBLvx9o4bqjCnRDdIvkHCv
kfbHYpqceWY1uMCm7fweLgvHZwe6rybOwTi+mr4gd93xImX5zGJXNhBj1xI91uLtnpDMWqEzKurN
2uaGyiTrydrDL4GKoFcf1cFMzoGT7nzkr3QIKZ5fC3UDOd1ClbnN26XZKK+rxpa/1sO3hn5VbeSt
4oiBMvrwIg+J5S/jTnE1KGUEh3Oor6l7/PFFq94cfeHe3c/z3zPpVEMOh9pWQWwaRPHKJSP0vn9X
h6aHQgDbQq+NVpG9juaQQISMdVKSkd7Y4G51890Jz8GKSE2tb4Y25LMmavhTAQWTZtgqe/lWTxnl
UAyDOJEi2S7GYyFvOPWUmGoXO5ZOwUKGQZhlD9XSOKkbNTXpjJCizATWHFvEeNoQDwsIVQrQGAm0
hUrPsYeqcG3vr9hHibzmIkxe+/gaNn4Z10Sc7xMsd2SFdN940V2T/LOkRUIF8A7D6mrfxL+jnSvV
Dr/sVBJEoyXgEus6ex2Tnta4hIaEeIwM0zH1xgXXS6ToQsSDMlWPdMw+LJk+I+BaU6mgT0iXP6cU
T1dv7Q0ucqflTf7jcPMVWcQOuI8KAJW+NCeBl/4rSXIxSPq/+E1LD5PT6r/ej0f0Z0e3GvczZTzQ
UHPdDeUb0vR1ldxHq5IdKNrLvs5Lw3xGE9FBDA07Fbj9ZDczR9b//Ep6G6svT6ddrghiiIA+Addm
jp8/8J+gq1qk/pcrrb0VNCu1EJkE4JO0BDyNY9MMCLd5uIazgIs5/5HK5BFzu5ZUPCNrcfhJfHmS
1RyFK+pO4TPxzTuRD9uzGDL2ZFk6D2TBiA1CWG8IwyzQRoVQ1KKoI3ueYCFtqgdVGVeXEDzvouQS
4qQ6NKeSel6HfTc1SbskQfVtdRh2VSzbufj1RXwx1ZvUEqibng3tdQZH4XLkNnUfUOCSDAkyQXGx
stmHFEiygC/iAyxMZEnYPGD1bem9PmGMf425E77K4yHassOtMhTQtG8Lau+7/9eDgIBSKCYPrBGT
QRwdrMZqKyIQywE/Jb3AdrtfYv1PPFs8wdVzec4b09T+/22yx2I6Wi9dPAnhzIyxJaJIJXzIB0Jr
TYYT5/J3QV3nX4IFqJuAB4vNVhJPyW11Xm3sVDAwGLS0t1vppLavajZoOzjo83InMp74+vVqYQf9
k5UPb8jmFvK2J18bB/svMWxxMkMuBDlTz6+WweqxAvdtkKcQageiahGgIxDy3NdTGmP35ENTXr+b
bzKRB1INbj96e6k162d8xKdZD+pL681qmP1y2laGg5wiNz3ea360IUXMxn5HgnkEGjN1HnjwU9TX
S7XIsjQTXGgSjYpnVz2AhkLaRptASUgf62Q30lpVx5yPyYwV+FRy+0IrFY8PQzQMzVguLnoMEFJf
/SNJnsPpCZbI33l5T0pK40bsdd44UOLlpqUAcy0bVU/Scc2tn/mPnmfFB3+yQKcvl4Y9TiZ62W0T
FjOWwA6LcOUGoziZMNGC541HGxdLiMjs2AZbP+LfydHMl9wUQC3jj18X2FoSNhtKozrtWhT1NcjB
bI4Awo50jkH45dVntZvMrP67bpqfzXPNS0dadlt+89aU2b6Jb90pZ0kTq3vjcV6JdvGE693igc7A
xMOKYSVrcYqHrHNVZ1aRHx86CLk0RvAsaCedOSh4sTByJXHVW9FtEz6+OiV1rwLn2tApa5WM2Sli
xoUgeGtOj+Kc9GGlRSPaYBOP8mJ0e+8q255L8KaGe8wXIpdQy/jkvQfk92yxLT1wAoJYSQJChkb1
/iMgfseP+6yitvd6HR0rQWdiiWOmTj/DYdBzlRjFbsiEBJMc45W/NS7JPvtVZwxzurCfqmXiZo5k
WHCMWyQcInhaE+HZEDjxRmY+WVeJrKchQJ0vMziZ9zGrUeI1YThzBhoanIUBWNL+eoLsNOCB3gCo
OThqFNtCAXUhb29KBmojyQdTNbE/TL6VHrApykUHDfkZVBaX+H+M61/iJhn7ZwVNMl7A0TUqO5qF
T+IVm2AR1+yQWv+evwQlHEDK72Zp7GhUlhFDs4+2oCmuEumLUdDGcROQ0FaZD8FJ3IS7gOppPpx9
q2dP3nt16N2yytDO6dNb/qwAM0t4C/elYHvvNcTnPPHs4EApXPQ1/Vi8FMZzMQn4GNQPJFjoUkGu
KiJe30RRDURsJXTQHmz0K7620ZqKUJEg0SzplcX89rB4SqnIbsL6zoJ2tT9YzFZBJ2YV0xat+a9k
53y4cV26BeU++MBQlmzNMshK7IWuiWGe75w4pU8dRMsaADAYiCMYOPNL8zLerCD7RCG5pMARh+GU
h0opD1/wNWwQhVhVtfYHbGbNxZ8ZEYc8J9mLe4PuKBVWMQNFmvuo9csVsoyV3hJN/T3Idzqa9ErF
InamEkJB0iDXo5wkyO8pGh8kEEa2MncFTascpGn/i1oQ4N7ENEYpE69yhjH38Fgdyr8y/yXiQXqI
7knwNV/S4FBj8YtGB7X+t0kQI4DyQuQc5wKMCWQ45l5w0mWViSfI7zG/RE6AFLqj5y2hyYIUQDMN
GaHAlaa6tKPICt4vpcPrR0xO4/tSJuZFMMd/EVNuWJo8Og5qs9ZPa9738t3ZTgSyldt0ogf2lzj/
xwDvaKftOj892C3OJZV7bFhN1PWiSKuZA0yZmdmi7wz9oPIDxsK8a9/ZgKVAIf7IApx/bQ7Iz/vu
Wxh4HcGjUSJoDMj2etJ6t01PGxTF8Zn2bBAST6wujbr865OOlmCT31yqCJASDXBBNZ0DlSKVwqTd
yH7Q2PxkSlU7JsRehW36INLCdBapoNxhYy9JHgDpcNpbY24ue0+jfBAGRV2bMMABKgXrKemAtZhU
qLX//CQq1Fd8axcd1dPj8fVm6ibiOJ/7XhP6ssVVHGkAUoGpPjI8kSoF6VqIl5emkTmh+6Lseey4
K5eQ/hvVoWGZzF6C6AzJ78PewG4kP1TLn/0RdQa1/s8w8IJbCGtlUp3O5vgEjIz9VHQjUnPw+28/
UGvf2zWb6vVGF6H5q0f/xfDOYxoXEZozX8m6QOc2X6hoIoFfNnmGIKjTwjF8hIBYLalWpbaLkqUu
kaYSwTZnfflygxpvLWZRvUXYHhEqSGjmm1/B9wSPyh4rN3RSuYNOZaZnZngTEbqJSuJTHut7Mc2D
K7O2Yc9UN3ATj+I8U+ZQzAQy4fEucIfiWvDBbzqybYVm6NEkJaUadyS2ewErmuchS1Byb+yx45iZ
Po9Tcj6Daxs3j3dxY+FT0LfsImt/6FXbYTn76V71jNMiv8e/pQpuUDKWaKOMjSvMG1UysbhDedqw
nEvbyjkEIA5Zz+lPEoJqwVgVzbDndhabbnZ8Pacl1cdFTU0cecWbRLOl6rn4j+VL2mW2s6wj7XOw
k6T0Mmn+MIm8hT7i4CKp4k+9fZmVI4MBXYpxhdorB7FeOccYvD4ZxryBcMhtM5EpbjnKMCq/twVX
cC9+4lIzWZHCqEeV/UyM4HMhuGRPPCMXD8nMcbaaFYWB+Pa/buHsjc1jGak92s0wZH4ZkumbPxbo
pQ0XVeGNU9WeJOPXEBaeQgvP0CZMqR384yAYsrWj9eDq6Oc8+sbhC9XdRjOIw4/2Mie5M0z9oynH
R5NmbfA/I8Mrgr1VmG3SLWRFS/SUFS4GIz3O9fRMVMD7A/gqPszchrb1iVQZ0Zhgtun7k1WU/2T+
ZZlm7ZLIxlsGzlxsxkbbGMXDhHRVHeaU7n6M5a24EwSbc1wkmHYOinFv5aKx5YTn87czM7NocGGM
2Gah50dHGfQXjS/0JFuToLkL9dXrDk3VdqbBHa1c/3dgGlYYAVy5EVbwc8332Or8fGf/8UiADlbw
8gGPHUb+ZslE4oCBte2J7euGtXsh6Y3VETrPDiHBpmE7gSMfMx0ldXzgJOgs9XDjMGFYTWIEuwPA
0Bn44MQ1iSclxYKVRVoqpbWwJ7Fz9+yAmpNoxzJG9L4EsCa0DxuUJLyoHZvcb9S6n3GnF+oLcpvc
/V+nNT+aQ1owz32m3k6dTleQCxHOjkfDR7842Ukle0GfGg6ny+rTQElttTDXz0mDHOfJrqbRGAtE
ZURiPXNMYoXYgjXwLbG16ARDuL+OLpUztchKO1HPIbAlFahMeaHhBuYCEB5FHR63n4c6daNUePwI
mRMce8nqzRu+CAWvPtMaGzXVOgIBiVAbP81ce3t9JmoglQKiXYl3e52Q09HaJV3SA88miFxVXiAu
OOV2Z7RRLbOlxFzJxARXnmvoO2DFrLdy5UjHw/Kor99sIb41z0ZbWh4BPMvZTA2eb5KbWk5oLI0Y
bIp7lKRO4C40TX/FglQfo1WMmwNpiAI09T4PFSIXaonCAAdMtU3aT25DMwhuB4krUACIGIXFdDmy
CbGsKTHfkoT3oez8TzmOyS65N8hDLFQ4YyYSBo8+VyQ6dbve+NvtwIedrXhonyFoGuuuiS5MRkTO
V40lBrRy37IPcbYXfW/nqTXQ90SUQXKeGdg1kzJz+V94p3i1Wxwwz0t9GaAOhDfIxXMLodXlys+r
ZBwRHhC2IuEq3B9avDf5vqA5OR5fJWc9X6GLVB4Anl5PiehN1NtN2AKOppw7O/C2vgQhagesHuNI
sIARRKsAQOp3ffTApKsYD1uZD9Sh1cQ/7Kq+ageMT1o33b38jLElbkF+uV1diZfN2vQbgRV2WmVJ
429Mm43w0OE5KCimF1nCUQOTg2KTy1w6+v9Hd3lHgJ91abnOn+3X7LRPFsYXH//61xB1SRwzaBEW
7VBj/9Oq8MCGJHIUVocbP11gzjXlDXV1MA7IfOH62dzQqbeFxYrtT5Lan9zTITPS5lYkVg4ZqFAK
5FGYf1joxXFWvUMtOPr6vJD3jVaMXzMkrKZEeiT9uNVIQg5GYbhUeSJkDEsR/a25tYBe2WWHdx/L
RObM4V/kMN7QVdgdVNpW9S+szE94sOGyTBTbEZM47/1OE5j8F1WKL2fwfzePmF5YblvxNQLgh6UU
LZlVZ7hVj6WFBywbfF6jXrTaMjy7zGoHjIh/oha7/V2tgLdo3cWyD4drJAB1eEOoxmcD5kAlDhbr
TvYImPWTV6bMDbkkRuVPtPplwMBfGQlfcGYNkyoMrjJENNPSukwZkfgqY+0fOnfVzevn+XSVcUP8
piWm0eq3wTTBOWTVFnMryoCsR6tU+8k91DpX3spp8TgQ7LlXsrjSiQU55nUBKOrp3Fypg+vBnsha
5QqsxviqGOGfDgFQofaov6L8hE4iWWPqER4UW9D72nxufFVQePlNwn6eH4rSruaFKRlNkhQ9zXbZ
SrxzbuKYf8uO3J58WG8POrCzBdX76jnbuO9it2IhCZ446fynN20p7cymoA/bNypTHput0mr0NzsQ
9pki6WCnyEg8gbzBrSeD+PWVonwbUMZaLSg02xdgfX8FVzv6W/mGbVDhGE3NT823SjW9q3N9DDor
FLYBvLQAfZyIHoCUdJuMWDYqMpUlb1yW3P3CAOzf00xjju08jBXbiMemJmfSfJiR+A5UNNMm4Bz2
LdQgo4JmTh4rlIk2V7MsiomJ9/Guj3pVFea3alkMzFLXb3mVzKmx0PdfnktHYAsz0f5v1CSCyq29
0zEsYt6WFWrdCr+ls35RCGA9yduv9nmdCer28A72+otb9rA/NYiH7c8crHN3jfpvI6VAvkOacZ5d
i1wMkpT2HTe51n+AomhgS83qgVPGqbcVe1oRLWygPIB6HfkZ5LqU/TFFObGRHajh7bxWSYoWhcOV
htQhaXkAXz0VOATlqWcmBvHYPbKx73FRDjKzhvKAkwJ4dMbgce7IwxIt/gKOgySxK+K2c8k/bwRk
nlY3dSGKRbbUmMNiScUyY3cmlUMC3vJMZ7nbB512ZnxhRszNkN4+UxKZ5myNwBcwsA6E0URYw6Kr
PqjLxsR3qWJ75Ss4yIRGBVkaIk0GOMrM7/l3zmBC1J+ZUloxk25PSMJ9dRyVBNGgvj1saN7hTbsM
U59QKSUhGXYUX1s/YgwsPx8FSdb/YwwzneZN6Ja/XHTNyZ9diPr5n80DLCR5cMJBf1its1Xy+XAe
pGLJnnbgzsHZsn2PzbSPQw5KRSUG4JJ6Z6Pp3ILIA+kJxtFNRJnnAZHmy0pO27J51wAtnY3La/Rt
R11kyg+MfEpuMnwudStwAGgv1nF+25oQHW6OYlXq2RuGqK4bHdKoN0frRayr2NzMroCK0ha4O2qP
i/TJGZic4a1ck7xS597wmLIg1v2E57/D5cFU8LkC4J0ssDeVTa99WYuRNzAx0hVWaMT5El1JENxo
KZtMuexx9EI0RWOPMboZW2g/ZgTAs7Tg0Nd7i8kQ9V1yWhOwUWdy29PT4kyICIvOYBiIAxIj5hMr
trOlMeKZDEUzr3McdDI3CZUGCjAKLQ8N4Eqve8unT8L9nwRDCAKnqEqqqRah5HtKbHuE86jGw/ky
W21SKE7YBMkHxquyg6pUYpjtLiUcv3N6RaXnk0MysTUs03X/RiLWLjMF64yjxgvAawKH2dMc2xdP
jqLZJjfaqjzDnky4RbX4PFTz5+T1W8ie9QD9/sTiRkC9tF1mSQhC2RK1zRpYVhoOfW3LtjteYHVw
l0HDv0cbBztxHgDRNd9J1ajtxHoWChBX2luQyX9vq2RQWdCACxEGnqAYstFrDK95YPsMIrTLZkYJ
Y8ak2ZsIfdG2Xq16iXU6LwZ6GwLjNNwGbgxxBWOm6YCUrZx2ASggnnyfFMi5qIXP1gppZfqbZyP8
631xiNF7vF5mGeFIQ8zdHNhdNTYS5RyfFXfuRZOXm98nUtOFV0ErhVHYNTif7tBUep0CbZEHpjFo
3CxBk8QikXASHK9xUbXLkJ1MVDE93Ptg0u1WayCoL9hshec31sM39oXcksSqBfgN1KJ+VNvFKkME
2e5ItomrgJ3EUWt4f6Zx62fmgFVAAWSfdvyJ28zlm48BE6nQy1dG7i26BLkUrvY8aB9Fe3LUsElj
DN5WAg4zld7VlXrKnsAkfe0DEDwVM1SGsC3ykzq5Ks0iVzC0OS9ysXn62J8OZQqiwWP8Wjr0tR84
Sh8DME5g3RY3tiFZL22RkNte+08g0wBB/6rhlDLQN6rClt0k7aIe78wgVN+ajAl/UbjbkJgeZ5Y9
iSu944OHoqGQvMOxjyYuKLLyJNoP3Jb+BMl0tf12y9I109KxkAcAZeTbKlJESsJK5tMaUKjZxiaY
zIkA7h6FuhsPoyud0l/ONq+t1B7383lWn3ab9NhZiwZi8XT5+tf2ZdGYR2+k7UOAaXrmqFO8XZ8V
M8To/BRo225Go/o+Y1akK4lQsb1+SdHn4xNcEMmtaKmZwd1T9qUNrdhzR49dL0kE4vLnsgMDWezr
r2Xutiypxgzi5Hwn59FrYkyHpyDKG3Yq7TBPIGv/5GDmulliAXxmztvs3l/7GJS4e7BRq5J7G8w2
kNFQGotd8fXuuoBk8v9W5gzswxzsotE/AFruugvVlKbXfj9YOI314/QlwmQu4ogCLoSizcJBHiUh
RuG/sMMmsX3Se9mO5o+hh0r/gs/DjSvmUODuBXPP10+31s+am/n5614IpKcMocnAR7+u20niC9FN
tPy5bITWLvnH7k2n/K3nYEVu10ifmocoE34cZ9YqynN4CDjkhqXJIjijAA1ftXKQF+8j5N2DuqSR
7QletShNn2kkTK/oE1Pk15rizsvyn3GcFSACVEWqUwT6n6IkvLwYM04p8tdB7/lvUoq+KhFzi5/5
aIenV819cb2lUzigPgtUJwmvqcQmp02gr3g4BW3ZCkqNc/Te7fLPlYssdvCm/wdjQ3dqQB3VGsKi
Z6FYcTJ1CAvqtWuc/GRCveh2FIQaCfqKCZSc04HievleWRooXaqF73+FcTLidef65aTwFvRlwWrK
UgTo/+YbdpzjkU550Hj2hDK6YKGoI/g/qWh47o3P/o6UeTrIi0VHnHrIZvL+0at3YJWUxTCzDzDR
+JjZkFdUfhT40kf0HcHyX3aUFVwHXqSyPOM+ByuYlWUTqngw/qcLMl94F09O4HKxFhrQ1t1xKC/e
GOjm9aC6/1ftogPPj/QjgFhyfFJPQGLWmR5+G2nFJuzKaUQmop4tpNF7KJhKSVBEtIW6qfcItpCv
sbBEDS4MZvF6V62AtxLWADNQyGQJa+sSOd289DWVPMzGyhMDNdhUfBpXjIYkzX/BIwQwLFTcH6IE
KQAwfriREgsFiQXNHziXZhHFTjlIjt1hn5G4hRRzVrZR5HH/u822aghT0g9HZVZc1ipyD24fAAiB
cxxLshv3uPzTrHfWnfD/FtOce4VZPvPR7iuKUDVrV95zuOeSMRfq7Zi7w3wQVo+kS33jKLnXZ5NS
FnytpacZZO6IALTFVRYTe/8ppYI02X6Bcl9NEdvQkKrCk7HVQTJYboJOdMeCreiPpmgV7PuEHiv8
IHGvydeokCAmnb77Py5ekjWAI6tVAInxZPdqUoiWsHgY+GCiQXahL6/qJuy42N9dzG3GtMOnBwJO
augd3/0VoGY/FT0PZZJjQxfHoEo+9bGnskcDLCl7bMEHOW0l/UTzUw1XpLPs8HoKhmk5kBF/obfc
ttjHFwHK+M5XRBOdK8UEYOUrz+LNXp3p+cLYMnnoA/p4aJcHcc/Jj5BbxM07mTdk+lfqNlfPGLZH
t4LE3Yk6T3MpeayV4MdwlRfP20fKFhGNkEyfW9U3qsk3XcWbbC9hrEhaZvmLzl++dasK7D0wTCHa
lzsOBXuJg20vt44Kosk0FqDB+jz/+2cwPHmIjFHG8c0rsrPa/u7aN6RUDhfMr5x89AQUvxvBgCNn
bgW/GjIM6hD7YvOkcK9udA3buNsBGXS7Gjl/Mx2l/+aCwptNAUkFgrFFj4psoAG+ab1Cuy59E05/
5ZepbTcFofQA4T8+vU3Pd0j/0Iy3eYh4aojdJbuv3kbjVxAhyYmhZ0CrPfLVbaCm++W1C4yupEys
AmI3L3uq/Ki2jP4zVC/9HpcAU4NRlrza3pD8iQVrJGGj0pUPbKNk8kKmUh2HjQ2JWe/e/2EQjTDt
4ZD2Dz6aGwGbH9CkmIh41IjxRYx02toG1QUD9+ExcDMV5ZxQS3Vj1NAavOre17VewNQPwgFHGtju
WlLLupPJrsu+2Sc1h7ePk+CuI4zINttgfv/fMKzXN71DYC1L3awQ3IpEzGOWU23twwW9bwGWLWHQ
CWkBRUrtA7VlEXlHMhQFdH98juxepaJvRgm2K8kK5cNvPmzSNZx0KOYuHCdvURNbmFGWIKnHASrY
emXRskk5abT8LIBFuvm405filKa6gEq2FQx4l+bsn0XXab9hsTSd9xKdno4SZteaEp/ofidBODNC
FXZEXjv4+b8PMbodrWGYRSTGIrZko4/v+JNGSRYzB8CB9djcBUst5MUnr7Fv2NKRxI1UyAFNXY36
j/+nkIOyoRzRmliSIw/WVfRv7ZjDDiqmIeFW7A2/7cU+VaHG7pUbXTxt9w04AvrctfRcObsHSN74
qlz2FBJGAGkZZq0oMTW64or28D2u1/vx+pslnm+s0fAf70Ufdgkmwrzd5Q9fpWSdWpIfNjENJjZq
L8aBaRsm05ADrBfBnjRzZm1TMXTibUx8PKpD66kg2T3zRoZtRC7fX2knNOk1fyRhvCHgPTf1vHAH
FobCiNDYLySApPUMym10fR8nu8eS98MpeIK3ICrX0uyiNGJwLVjCH84Oa/IH5U365c+jkvikFdfv
YqhqbaR703E+1eRfdFxgI+BZDNtNxhRE51EHaLgHKoz0gVXIa715fd/FoVgZ2VaLX6Em0+bU1/rL
kljwX3dXgQpY95VayGyIAPdvsNgQWFVNGFDyPXct4TvGuSbj1sSYRFuZKKsIvdnjXDccQ54Ru1i0
vkoVOprttRUBLpalMuXMt1GO0HLST4ceW7i569tXqJ70XvDAmKgR68fmvsN0cJRZJEt68AxmgCa3
ms2N++TyMnFt4eEjM6d36dvzRa9ltdwSxOPqZ43bqnprjO5wNTI0DC/ciIF5ht0iB7NqqCsCj1js
ecPGl24ow+rdMDe6HnApBlB0txPLxja07SvfJqa+AndGuqfAzVhJ8fEAgPXci0w1xt8SCooSspYb
ACVJGBWQNdtG/+NTPCc+8JzcmTxW68nfRi1HCjisQFTUaUuA8K78mHsHuGsx9znPCIEBvhAwpTPq
/YdrI8/5/QjQobe+rib9ad5AIzM0p7549PNVVdrXgtk0+XC8O0ssU48R6a1UoHBi7ohZZWpZLg8y
XKX58v2jJwL7/64/4bwGxjZ+A8cBoETLaY6O54fqooZZGOZRu6QXcG4pCYIov1++uH0tDSvJYpvV
aK/k+VHFCqzsehVrDUz31GPgWaPU7hvJcQsHaVvGH8yMHKTjHei20S0W44xr624O9/74vlLg69s/
fjTXmNY9GihjY2jbe/FTWpjiaEtep+t/dwde0HDHuSOIGr/wcLYKSFQMyXmUCifV23ZK2SBBZyxy
gekougiXPU9ErfUUX8CwN+U1bnTLBqgOXpCe//Gh088l9pibrbfc2NzVjI6qEV11p3YzvfqmDuaW
+wQOlqJfkx/dezam1Fnc7HpqrJm9IaZYf1XW6aeN4GLazYm2K2/NYQrWJiRuHvzQUl+w9rQICLZo
4Wbqy9Q3qhP2wyaczfSxTsX5nZcuw/XJGGr9GX32HjCdg0fNKNDWJO1sZ2/Tgx1QuzhbwIgYgw4y
2zaznQNPQdgJZ5DjNPhKtEwRKm0y5DFeDX4FZX+4D0i6j/MoW4JwI9MV0EAbbmC2unl18jjkLVvQ
SQuH3lFAmZY4kZkG9s3E4y5zV19nUG3Al6UOjBKLMJV+qKniVpf4waKqYSnI1MlCd0DdDtXW0xKR
VRDy3DoaXHE1UB3YhicaF20f9n79cgCiI7XhPgMTJJjcC0WB01OUJhC0LBeYyAfv7bNXmk8AfpaG
ZiAZbRT6Xz7HtPoEFe07kYoKsOy58aaGFphupBoWWwGlrLod5cNex6D5NrXF6Xen6Md/DJVwS6hM
gV3hq/1n+kEH1IG8bTJBA8cMgaaeVDsrBDbgFsjSPJHHUKA1yUFeNPV3pAxQQPCN0yihzM0GczQf
PvL5mJrS3fBbWFO4VwGu8WehGm9fIdpGLhEcNPc7j+SqdkEIzexR+JPnF82UZyZz7u1oTdZFd0Rs
HO2TOazn6l5LWYWy2f1UHvRgsKmhZRc4Jquob/hbx8TmmCSofYPJ7xKCHGT+61IiSUXOfnNfp8r3
YMNAo6coYbzMyi7ysoDYrFHF9F0YXhrcqdoEu4lZ9Gr+iX2ikd5Z1q9VEh8m41u6hb2FvRSehZ0H
kTwHZgktgmZVoGDkbhl4p074A2BvxgaK6NGdGaAUPMh50QTnGabC+b7fVsn0Y6ubh9msD9mFumya
d5XyktvVn3DL/yx41W6eXqL0F8l7tEc7tiAqlxS/l23PmH6dGM6fO11RpBErMU7ApQ8SIyQlv4RM
Nc92+NFGzxdXFWfHflXdZTh7nb0KwsYXpblJzt1QsZHcWWzj1aX/5eLwYRLNUEM1fnf7xVqKHjJx
FPgUDGSDgO7aeRprI2cf54NZPrJmZ1gI2d5nBxPASjuk+tgDbaNdYfvwGYRD303T7RKv1YFb1FHN
jCFz+JozhjOMcoqvVkp8bui7G+eiBXqXo6ikKXvwT6LYbQcH25pWpDRAAkm3uNCwOETZoGXx5oKB
FQPU/tmvYOZtZ3TEIQmBZBg2udjjt6ZKlzYJ4ON2ORXaSgeLlVh4ay3pw0BDrwT8Th3lITBiJuli
Ppwz580dQDTRRlDfF5U+FLeaBCV2Xnb9CmQy46Sqsv1R5dRwsGA20TPq0v/QUi1YInoRykhafUR6
rg941NCcg2kgo40GY/sdgpXSPe/OBh0n1ZrepcqWUgYQ1Szi526S5u72HVbIsg/8s5TVuKRxTqYD
9a77hH0DwAfRg2w04lVfj1W+mO1JZSCpCUdtHnWXKgsutDaSr7JKqm3Lm8CL36H0vr1WCvDidr9d
gZIWSe7jLKzWgKv4rGRIwumaPG0mM+/JdhRU8xGLAiG1Fouvuxj/S+qRJXkhdRj6gtQJaespMxny
KHSu6oZN+ib/pK7elHNP2J9tgZKZ9qXezEQ0CohEv08tiuPVQEOotkBxF0PDKKXyowGWBSg6plRl
Z2l3Qwb2+cX8swo79FbmroyM2U34I10ns5jXGTvdRWMNUMKge9Xq1GyxXmogYa3rbBDE05gJJpeE
4AqbEmVD1U6a+SbKcU2S+9UWqAlfsOlMEQPVwJ/pX32D4fDUZf/e2P8ZdAq4SZ8/RCDakZzFhUnR
cP57NZC3WRWNn/dQDVt3q4eeX2eLXp0MAI9Ubx5I7L8kqn3rOmwESNnOUMG059xOp/0mp3j4gtm+
VkmEUhdhHSe8a5c9Tgh8gK31LcaPrYvK14zRZUJrWet6stF4OgJrmCIYrQkZChIONL43wvb5xH75
7732aJaxv+SdoBIfJvabfF5cFaS7i+hVjfu3ByjLQaIYpVjeGxbKZ/XI6ZqE4GCGNkHT0CmE7cJe
oABuP+zjxcSwVy3hJr18fT238j1ImOX4NLPxHOfh6tvR4wAS532/vEg3rUozOHa/8+ZeEzS6t7+M
UahWS+xdkyiEln4F2hQAkGA+7HEdloxELYSUvnyNHppE1xpN2PYK8xPHYPTkF8BosaWuVJlK1gLg
9nKY7VRF2pBxzhw8lfiCzBlGlbp04rK2ePEm7M5t32fHj1MtEHnXXOPTUDpQJumUXbQ/owNs3UWI
O0gfK0QTV5rYYFlqmLkxq+CVMEeQFLMRVd8lihYujOgHiTxbqXzDOas8IkGbpO9G0Z4rRvXaOHK0
fZzPK4Is+vczVis+Z5z/ccbTEVQ9Gmbgkelpo8OpjLE6rc7dhfDIqpQy5jiA6wF2zCIILg8jiUlR
dxZJcGSGT/5D9tzv/OuNLfVyntTutCwpxmSYAw01SpHqu0b28WkSpacs6+msawRb3cBpDA76x1W2
wOGW6RUCy2i9hImn/nJSpNMAgGSZl1mYGIxCRRoWlEwnD/kfaCPWwUWkDHo2I3jrcLDgGwBpt9Be
nDKiMlNSJRUwIj8LT5LVWNrPOj3aH95GOGNERNONSSmU/dP6iRq8ip8y/N4LiPGNB1SE41mkYDes
eeHS9D3bMkJf6RhzLMDhXuVy7rJX2eFUt/gBlNNDQDrID4gmMgVj6d1xYKQKQyYLdxZgC4YMxUgV
IhzcIQ1YQF0dEheRO6G0sjTmTsTo+71xYXfj2nTqTfV7UTjy5EyJ2Cb2g0hchrDqvctPveQsDABR
uHFsfHzFQiIV87Ke1ymXcTjM91qNsLKRoboCH3H6NkW/qvtwB7OMMrjr9GG2gLWX7g5F8A/zzipW
Ner/6r9/FE4l6KmoH3JBS4qJzGq//NQ8D7TqfijYSbV8/TZpmcwKl6qfhhfQ/1dN9H00dNoyod1z
2CrDEMwT6sntHf4sLWwjiXHbrEBGKTQfYB5tRr7MSclf4jfXJE8fMgUJe3QoD31Q5u9KpgzDllee
8q09/BynZ4xjESxjp3jNnxHG8pcGe3S6Y8T+V6NrVIYk1qlOBf9NJeadGyyMomAf0Ivphd0pGBWK
EWZAk1dHzaHe0LiKvA+VFdpx9CfVMtAvui3qZ1pHrYO98VPJv8xHIWpDUMHr826NIMoi78eVGB3v
HSY8EBNZCQi/i0Wf4oouL8/MCJ9lXPebZR8zT6NzNO4Bj0G2BjyyhJtyFWPAKnUlk0+5IcPj6T9L
hLooHN4qkKpjOJgEuqtyVDyQ5Bkdfd1SKPfl0aFq95VoVMZqgY2q6UrRTaJDjmypyk2tgQ7HM+bd
zki+edGE1w7aVVMfWHK/2YNigwEG5jucpsLeOO1+vG+GzJc98ySFb/WGI1JbRodJVT11hMLdVVSh
1cGnFrOTyJMMXbDx6S1tK5yxDxKJQvfz1ix2M/OuGDrYH2Jr0uzCMDZ04aQnIfarm3QKGT1y9aVb
hKCdIUFWRP4Fy1aOPkTaZ5w6ktUBOTbQ6QN/noL4fYtkm4QCy09PSa5g7jABbSuFWqw0aIobnvlN
F74+xtNzSLr9mOVQevhJ1R01DL/PEmun/1KENPvQFFMrem/ELBTDxyLHf/9AMXJqJ8ueTpIh+MTS
JYditpKEhtSylmZDiAzbg9fV2RElY9GiGhg/m8TLtvmgNFdlAE51AI5foHEW2mQDRdwaG4QC1jvX
viKkpCfUsTGS+NFhEWq1dnVxOYIDAwSbBDoLwZ+sM8Sif4hEBfmlKgCZftKdMLi+9taftjed5Ez2
e7bA6l9hPF2/lVsZPxtvl5TrViQUFVCJ0KJEES69n97kyeDM6aomD56lEyTWA/kabGSaU8XjH9mq
g/tRNiZrx2H0hqdQBi67l0hS0XG+lfX5B8sZmPi0jKrY8j9BpB61k2EpNoTMCaeh+RQGRWlK62rv
ogwoL6SYY6TP9bTfoCIOqzor4mzD6cSgMGLil9JSfZ4cx0GYNIfQzv+EbfqFE5cFrLvOqoXdF/Oi
iXbAz5Vf9xy/q/Hnayj4TLLOkBwqe5+i2JO7/PhWMKfL+I1SVbQemu9DCEJ768Nr1rpDGzofdsqS
kx5w1TklIP6okY+P22Yq1x71OEq5kkLaVPLJFS2dzHdhpORkLQQ3tYKS0ZTlGDZ2sYqx8zWfDykh
NqMcE0cpPBMLocndbsRiGJcspAOzbMXPp0xHcO8FcOrW7FSmvV9JcNbdniVy8BdbOtwgMQaCBW8v
mAakAB/Ugu2h84nLCR5s1kNkUMhFtnC4Z1XjYhZc5T9YbavrudPA4SNGVFiXm9JlMoLLECqD0NLJ
fQ+i5GLCLRNBD2oyURpYqDADpIdTDoDFnJPO6PictmykhS7L4SyTkwB1Dn+pfpb4JmL0gDv40vQq
spKNFdrtBUaYi05iWMmApTqZPPaycI/p4DjmJ12pG4jBGY3w8vFgTsErCriZkyO3wLNf37JyMoM+
7Z43lTIsePwv7op+Xw0gbYwkzQOiGEXgIJkTvpmN4/+WKqTJgxDAWVhhMUWQ9uPaNLDluFnDHCmJ
jo1CsPnP/m6fnRXdDITCg+h4SWblALphbyxfcMprRk6HO4Vbd9hDnZ02C1a3HMR0pUXv0H3nk7Hh
MFfp4SwzJzvggm5o/HuVo5pSkSbMPqXLYE/462JrHR1kMWYvtyswKbdJV0b4xz8MDrHlZQgnyU08
qLKa8dKQWXJzRUlYfDKtxb9tNB8rhGmvJFtkDE+Skqwmz7pcNKtVBH+r0XrBy5kNu07C3dg1k9/K
u5n4X17IF9/VQax0Bu4db8Wln3+rM/rCH2EIVmxTpKwhTsgHG4KBo9zUQuNXnDib16u996mO8oWM
LqAY+k6Kx9+H5IGGSUBQ0nZiUEiUYIUHtPyaFrqNXX+V+L8eP9dTQtVpc67lUxFBX4zhwGJuXxgE
deJpZ9ToNUQdEDOsVcIreIxQOfubjfSq4xYLoAOwZ8RF37URtpamIWA/U3IK6VBhwdbgFJiJEQVa
mbDbd7x6iK47Ii7YC8hWUJD/oePmnwDm0PrGc8vwNd99CfRwHacUcz0P9YzEREDGK6cgnqdf2d+1
HfnNbDj9dO6Ulm54abxO47B4iDULJzx6qT1M72r+h4ATHxP4jN98F2hbg37sHk6I6Q2HKzP+mod5
uXJuhkTrz/qzZqAMMbBLhSljt4KVR6XKQJDz6o4d2Zcf3RsX/1f152s3EEl9YP6XblLfut55MI1Q
2RCgl/ayyEntL4vXem2l7lJhYCuwe4JVwF3tNJjbX6Df2hJ9W4s/JC91VXWO4acPV4lqqtb44r8s
D3LqetKjR+EE1AqlHRiz90zNcCVTSzF1WVREc3LM4VzYiYSnYpu909YIwi4SDytO+UtN84DFdu99
M1OFywQpcyuP9+/hpk59dtX4jZfipRPqMlQ71bgYPGwA5qHv4ylVYWzAkMkcnuWQHDWjz+RPMkIF
Zi2PhLI5PlIzsPZqSmJPW6gHg795vYF9lHQKII/mr8PNy1JM5eK7tWJ1gpawN3zLU4kL4toNFutT
ufXUCnYz8UoMotO19LzdRca1Xiyy2TGd+Yd2wyW+Gvn8KTndk9YKMU2xwqzXfqTrTqwk8aGjBnYG
qDpk/rqBPT9KBVmQk1BmzbDe3VLYt7xgnYvfoJGqqtyjXpBOSlsWFUtlqmhaA32HPRTA3J/WkCD4
NxLOZ7kJZLhFwoffPQk2/TJbI8rMH4eD3JUPCmHYR8SPQPlXvRWdy+n0EZq+oFS6uLePemYz85Rk
L4RHJpWxkVAojnIPP0PfEY69zWZLKUl6g7+QuCT4XVecaY+IU6lsw8o8z8jWY0ezCNxYU+gwn+rn
Ok+BDZyLNYjg6FPyr5Bj4A/TMqGvQ+x5wycpzWe8vTPzVY1YNBbPvYRMiwGBLgy+6EzcYkONzUZH
6vVPiVkyZ1fU8s3YEyHC1JjsJ46cM7E22Hrorg4znqp5pD6BEWVvYS01B0nyNCFAFcvie7ARxAXR
atHCm9OCyPo2H/T2d8/97NAipTut9a6ugpyRvpfYasTr2xoJHlXY3PsOFFniuxHhVBS6BckjPkvr
8XsJ6s9fgb26V16tQ42egDRGhrFf+UWpj4Z+T2j2vgnlOqohFGAfO0/kDiTnlmJrxs7fRXUrnc0c
1uqcMc+/2FzrvW0YfQQICM17XCaVzT/WCamc5udA0JoR329EG0LVVFeuhtb7EkzYJf3vvCyvlo5o
r8ePHLrhnoTu3+C2gBM5gz/w1AdUVU4iICegEuepDtxplc3MWBVDR4F1ujQTxk2V9lSP8QPpGhH9
MtQPhAUVH/ui0w9P7HcCUc4Ma2RwATa5odkwd6LvvPUvrusD7x4rYUNrN8EBSOpBp1K948DtkCjH
qnNT6QGm2sAwNV9NwiV0ST0dZyAI5/Fu4C4vsyhDY3CJV/ukv7azkrnLC7fz+0Zk3ITXxnvwtuv8
HYZNxKmRzKo6U1viHnWtBtgOpFFHxcRo2Wc525fQr+QihNzcLfLOdhJZYMDHBW8FsyygKJpaR8HR
fSHTMg1HXhodahxCPz+h1rn4gV6WFJmm8/YPz1Ph/n3TuS0Hgo8jBsTKxRW0UXY/qripseqWhfsN
+KOaGHeRML0jPTqa7WoeU3IMglhNivS4pRqpL3StIQuNrPFZdVw31U92RS+bhrmtg3CTbPLddWS9
ihl0nU7h7rNeCJPeCd15G9/7GLGmFpi3NAcfTyvJ89LSqy9lr9vWVnbtEBD+AlTCBWx/bUjJ4oQH
47f08OIzBe4XzliHfAx7vZOaUXjJMj+qcu7sI41lfNJwRb1A5f2yW5E3DhCC3UXmbpTBfMcxmF7H
GBEDF6GqgG3Wi/qU9AjrDCMc/vpSo6lzdQkiPuyfg5jEJojYGEcQ5qk51J3vS1AhRVjCNcvaeGWt
lEKqJqg9p/xw5E4U8r7L4UebHYVJ2UQUebJLp39cYD7xkmgts7fgJ1VeKQfyr3iGdDdMPgUAhNRf
vlzkpWyLHXE6DmZvV6Y+qf0ZdGNziZJBfkQFGvvg3Ip00ucNYxJzeG9mx3pTJRquegn+z9PSFoxp
FFungUlCnFeTLX/hx4y/H9OJb81g4AUGtGWfeUsxQmevPeuy2XU7xc2UuxwuJDbjUy4NYzJWKGAw
BWiU4M3gW70TaybdYig0rHtqSfJw5KDlGDH5BDjcriXeIuxg1xah0xn5VZoD0vA++2iYWq22sI6C
iYZ59iy2uqIDOZotexuEHIjuSl29wb0UzigTDlnj/qZwlc2H3kqo9lSQDjb2jVqFtzXJdHgHXmfU
ukK6PD/tfzRaSscV/wyLdWjLFWxzgQyXp10FMDXheeKvehldl6tC3rnmjfVxCZLGzdnhQNF2emPu
t/6A4k/Ke+DsEaItUHkcWDjkqT1AzljZ6fDbg/ltcZEbF9Nl55vTNpkZcV6C4q1+YMxqbYBmrOiV
WjFviksZHiC+1PUR8Bu5zazsxVZl6PANAa/oTkFRFCLfcKVUwoHaqJRcA5TFdr4kPKJo4DcZMfSN
RZFd5JBqLWASjXtoIcEOBYaGJ6TO8DUDD/k+YojqQiZeVBZ/LYgtUFvHnXF2wfjiKMgSq4AbfXq7
/zO3l9pDhmcy2FRMniT+xIym2xb7LnnXh4mQlFdTBwAWf3yeLV1AlEEwQF8fLIThyMojucYxvFZJ
sArNxURtKnJpHH1FczOIlK1JmNPr/76NNo32Me/G2cYGxty1q2Z6Gt0363hHCoKC8MnUcxZpJTjG
y+fVrZD1Wbsn5ZdmCcRQ52xJXF6RrnZwvQaF2o/6xgjDSLbDZ6x5p4fDlxZD1jG9TdfBhXcJVIYo
P7qQ2JpmlD6I0rA7S4oybcoJ+X4KppBb2PmY67zP3x6wq+NbnHrIa+DkQ4Tbs93eDnMBsL9poh5C
X7cQLK+yScmlR4oYHIRsy5nxjx8pwwjvs3fxfX/e+G5SdTw0feEVV9enPX51W4ocBGi0Hen+gsf8
V4ek36BQIpZtMq+auzier0t8KwdjEYqoHyF/slCARPPOWvcIAvK/Ze53UKMUi3lIu//XzrKQr58U
bz1IlgMnbdD5v876QseC1xO6osnajuCgIh1PedJhdbNvzBb5K+yv53nPZ24pDEtdLMgr8aab36oZ
2HecBnaEzDhsbYcnvG2P4Q+5FOjJp0RrJYSG7X6sSYY7V4CQ7hhrJdlo1UrODsnJoUVsqzt2G97i
i1DkxGrSseV2+hFbZ4DJqtfuJe/VfAdzjiULvFL0H+vQBXCQGP9hyFDjQ+caCniuXFgOc7Ueo9X9
sbmKrXvCx189XiHQzM1JdBD/krFCfP/7tcb4mI5QdMqblpxgB8EJX4QO69Uz5IYOl3d4l3q2Xhgd
ZF+Gi4UViv+AEBr8LKxZ95Rv746K4nJuDCTa9D0s9iI2iY2deTRaBNMR0yjAJc/hnLCbF+dxA+gv
SGhb9tKNfowWB7fd33MtfJyC1w33XV64oBI+7r2v2Ssrw2d3hJB7ri3hyKKwSfgwL738lyK9+C/w
KzFEm+4JsdsV/SeNGDlNftpvUColAbIUEZYFnrdl/+a36cWUgvowqA1lSCJYGne0F9dQWVnWW2dr
pOxBzSYdfP1Y8Xdzd26lKAINV9MXfYDlqHNHrW6rMV/QXakwaPhaL0a1BV9YEAcdJYJaE0cNdbkC
TXo1lJThWCk8WBxMnzDUqiFn2w3Z461bhbuogX18WUAI1LhC1z2dDRHpbUxHOWjp+7/VhLx8eMQv
v6bg8pooTbL9jTvsYRyEOzAgausMqZX/PYpQf+R+coL8CAtlmOFLEMOk7WMOmZvjYv6Tp76BMYpp
BX/B0qWWZM6U4BSUCKSwvh5Q5ZuWsFKf3L5Ay3rtCPNtcIaXjqygfJHOosdOa1il7k0hqFChTeDt
yifI14JWAsW11zHH8cyTU6/61rE4h7Bn7lIypRxCelhPRrI26skItrJVV6s8LEZyAe/8n4z5qaoT
TEoFtyp/aGntphjyff9zXIT7adTO4XWaPV7zSHkt5i8wCecgjTbEAqaCBa8huiIBnkrk9+yI5wIo
bgLmeUqE8pMmA8pOjAWhrb2uYtkMYZGv+XCrVLTX0IDc0qt8VOdl5W3lEKNmKVAavohzgBghLDdn
hBttY2/W8EArigaKzvYiOPsSrJLaBej9FnJkFR/GJsjfEpvimfqmBDGFlGea4+g6Z+FA7RA1wxOQ
zd0qLhVgGvuQWESnMco4/EBQ7z8GA+mpyTB52Nr3tYq8FTGh7OoWS798Sd9OpfPVpFb+TkhQR0k/
DfiWs2/XkP9ej62bSWgXLAMkFh8QBwDMD7i548ET7RQ6fhB9KDh8jJirWZ8r8gcVocr6+DvqrxWU
4zRYUaPHj5KzzBrxzliwyTJm44GCTlJHQKpyOShqk8juZOe3NRIvzs3hub4/NmnL2CK/HopL7JCx
SuryFCImj81QjyR/5KHEIxVOXWj2w57mY3RkTL8+9HUo5D+kgc70KnT4nsDwpFNfrjyJ7qrYXou4
JLngDYgyU1dywaF3VvWfj7iSvNDd3EJGRC7lF0BOpkRryTDeYf+tOcV8p4DqTI6YIf2BE0gDnkd2
wsI8SY7W12BEyYow8S2MOkFA4dvIaWw5o9dgQpz7BGz1rLmm8N3YSeweNHgOMAxVENGNc54DhSgU
tHxCkA1YDxmJE2t1TEMNe3A1tit4Vuygo3/TF2hjlVg4jYIIZexjdhGHMjiz4lLvPaLDr4v8bCJ+
JKENcN6Hju58c4EMuIE3Vxs+buSzVDGYsv6kcvB4nIWWhjf7084a3mdkRrcNCnJM5Q4enRhb/fSh
I1H1nETvJotHUbxUlHLU0lDdggQAdDk4QJUwwStppSdXvBygORxQrs6LUrG9C44TG+KFKUsnYh3v
Bp9/yj0/Pcx/wkqth/MV1l1m2rw/PHRdfJqP8ow0r6PmGjkyXkut228a3O+Gh/ziYQlw3vrZc7gs
r11V3V/BLIMBy3onlNtBRdOd4+Pc5smKCSqEmTPYCpo82ohwAW9H+yvyv9F0IvJep8sOJIA4e7Un
YmOTgDI6xm094rlwGAEgJ2xO30z/HHSaOoG7hSCMBw7np4s8OUO5VB7n45jzZhI/cMszfYrXXys6
+TbkVTdz6qvVr5Q27eBriec8GWe3Dx0VGMVLThmpfUERXsuYBcT/DicaNPYaxNQkNJrKxQY1wCr7
57Z+SjpVYFYhQq3fpkIJxlClMy0QrxVh/ImcZSDCd2Kwn5c6/NeBu6qOkg7vDc9Vga8rWySjTN+M
NqlFUuJzOGT76qicBQboiwEElzJS/w+wVnMAvXRH+OKFRvdnEuU36+x+VRGIT84AF/bHmR5kRabL
Ny6/HOuI4CwzQ+klMiKrSucaIRGyH3JvNsU04degWuxPmfy6VdouSqxe52UCjbRN5Y2qrnyAAR1Z
fRVTUOyrPrWqhUfdRYFpAi+7j8PVwrSrX7H6QV/UA+yN57Mu3Or15YE4HI3GS4F1IK1HSwj29Rur
RD4dxxX8jkwMp6GLAkNVXhpp36C5bU6ehqpw+EmBEtTQaL3bHjQy+IwRAkEVheIXXkpDhgyX10+g
1H0myaomXkZhCY643kY1jtRLX+ARbOZuCsN5NgqzSyipipkQSJh8UtpVYKP4DlFZv9WNFD6/Ygx8
SXm+6iMKIhpuiGQxd4LzWm3RRZxuGYmnDfWwyMFKdfT9eOcqkeMoAxN1oSbG3AQ5+1+0qiyzyPOj
IbGRZFZYGE5/PUVWgpoTNquMcSS1OkccHNnyFdkat08VMK5FulfOQghwIMsRAEW+7X7CyXY9+c0c
Buuquzn7V2aHr9mcRkkCEJfJZbcUkMGREKe6D0meIRF9LWyJL4KDM6cX5T0GHEC6eqABplzoVvrX
qhhuzgwClhnQq6ksSltSENU/kVUAVAR+nXZndzZdsLSTX0bXRlJcTn6zavk4b6gCMIDJcqspZHeO
G3yYp9IW5CfBVqXskNmjOps0mUShzRo+oiSEWKmYjoPqS5Gih4Wme7SUEgZ5e8OhKouXQqFj67qZ
jFpbU9+EZVbOyRGglEfe9kkz/ONU0wseIX/W24iku3gIgCRtJz0fx3/orI9xxeSBFlwJC3zY8J85
DY5g6lQQl+xNgXqLyFlGPMZ7ohRforTY4qRmRHQsnnYFRZAld5J5y2uu2ir2B6ZTMoo+/5tjJkIS
VTWeYMpUOhmm71NYeWn9gZLm8qZ+z3TqKJtu6y5lu88Y8j7wju3wkXLS8C4jNa9ZOq12W9e8ll4u
POykqt+UQuvack7ExLC3rUiWqpSVGUBGRgHPTzTZpzcLFM5e7elk5fA/S2kXRdl6gRYKAs9Kekyq
UsSGhOxJIdeIFeLNWA4pZX/WnyTPKOF5tJ1SRtqFAIriYx7rXm512aDwOvj1xGPmLmvQE/zgJgb1
94JrAAZe8n8DVXdxdIDiarbSusi99qeD5Ypxoc0heoO/N/sdrSXgLy7jH4uXuyN/h4dXkNmKTR2X
w1lJJ5LfsloNvIBvoiafhkn7ZfdSh1/zzLxeJf2rxpVoKzsqKLKb4G8ZM54i0prtV/a9IoZaUwdX
D7dcWub/kwXIgEdwBib1N3IhDAwXqixfoN0LtptvtRb0nICJk2ZhKEQs3QKciQEIS0GfxcHglqcO
DLprV82G/yTUFK7P4/5pWsylv80ZXDg1d4OZu/7kDPsDDVe/pyV3hLReO1OmQS8Wj8qaK8njs2+d
sKxRsFwkV8nxqgPp8L1d3oOJcvH4Uo8gwbARn/9RigzvsjaiqUMxXRIj9IKTzR7XQGgAh/tqush2
39qwPseZLfBPeeMPYxU/MLfm7m6EAIHThEVZIoyl6SYeYJUJWuTHWgTAoE4Lid5TRlD3bVuaks4s
2BQbTk2GzEL6tYXMQnzR5IbPFwdOdd7pOoFRn7MlyeYnLRNBiZ8dNuTHALby7yIYYnCQbSoJrH1H
L3/E1l0EE/LoFWm0H6f8ZD3SphUPkDGLNCxYrqqRFiX1ixCpGie1AFBmjM4+1ifFJGTNf0Rqqpz1
u6mCN6l3SMqbQ7Yq+FEvBtsc2NM8JSwEPpKMtQLH0T5OGOOjiNqg/ZFnGvP766WkG4UlfpTD+0fF
PHyfxUM4koaMVKdiIa1skjO4W43Q6YA3MTR+jCOLsGx+FGjaVQhYhcZxbFdnSMmP/0Nt4S2p69vc
VH/AtXVHqusqr7nSUkIE4HFeaUw+8IRyR5DQqB/JTphnSyCmhZWO6qDEzl90WJTmfHAHBl4VbhUf
m/UoX5R5GHMuyqZJE7wNYQsZd/b8/Pl7YdvtDntOLkyTX82uo0ENcWi7fOIdrBQUTUHc0cVdrNxZ
3gAVtDqRGI6p+JV/sGqpwb8bQvYWJiAAbXnCoOUPQgB4AV9u/1xn2wNGZEJxM+AXslArlRBr92Th
teMmgNcC68emTre0k+HAkNcFAhbBB/Onf950rIKufRTICt4A3p8tKE9m7BVqT99sPNWCHIZ+E9Gf
DaZi4IKEDPp7B5oUx0Qg7ErEPw0wG27SYH0QNinfgb+HQCnovTggX0U3Y1xUa6of1lIrhTlkt1h6
PklMxvzz/kjL0yu04nsKYwzAjPpxmIxW8TiXNsuYDcyh+ZTGisIwvxrOp7YPajUvnifuljRuf5Z5
+J//iNifI83zZre9l8fQy2wD8D9Ot+AJTvOYyh/uGTdc2z8ZRzZ2d+3tDTocE1w3AgFkCU5+EnPC
zeB2W93oy/Jxb+xOHPjwCx85dW0xaH0Vx1jD8unQO+brYTxLGPcqTMgzxjgNuAx7Wsmv8JnPx76e
qJmwLpNwLEwxISPyuhaYlgU8Ivb9FpG0iwQN5FTWUc24hvsMmYUGOLPDiHsddpJTxHBh2U3gWuwP
Ur0CtoBRSR5SFgvjXTOJpsdtWmhHEmpfVOwQNmxKzLlgnv3Prg3y4bdF1oJHWbfN/jqM4ZfTQUZz
QAuCDYVbIwFod4gyELH6l6hC0mDgZENjpnI/Ikr1qPJ2vyLQU6FWTiBQRZaHKUxzdg+0rToP7AOp
k5wnw9+uuyTjWMjh5UDgYHsCWcJ7FgUu44at3Et3PjkAKghq93my1aE5Lp2ITR/lHPLzfEOKUm0k
LbI0CxTyujiit4s7J9O0eS3cXt3kry6suAVxD6bDrhk5+lsPxkN8e0HUHOfjvtp++K2SKHV/btUb
S3W7uuy6Goojsm5VtmlixA7irY/h0sMnbwT2VUQcin7pmlbdGLnB0BfZKxgktB1wHbfKRr4JuR02
OCy31GjNRL+aZESpGhP/EnPE6M7qVvDWeVl1mDzzoJ/zRxlB5qHg67U5MzR6ZzxLNo9wqm7ixDHs
24VcZRhYBPXaG6BFgNZr7Qw3Z2MRi0HPTe4YzVVlhkXHZys3KjloJhSc56aZd/qq/0cqjAiawxY0
4gZKDfwUFOJebgCzwoGw4c9S5NLdncMMF0TAUlfDS33UlZ2U0wlbmOnQ9e1EF2aJJI2Vzi9yVkh9
xAg3C2SvU2ydWBdeMv3liYNmATIuf2MUmXJXRwbNfAksQYDmD8PWwm2osM2a1u3OQy8i1XpgyPop
QGXfFqdSB+XDSMVZecsIaciKnvYcIuwEnsCPtnf0W/vbNnXzOARgaPqwVGrflDTmMQbB1tdLXa7p
56aAfWoxBHCRU7/YmBqsV/8/aIfOmFbAx9YZZbBX0w/BR+hzHeoEvIE5edTpY7oncesn/wgYEWDx
eS0BdmdW0K5ohmr+BoeC0TJj5lo+Q98DVg9caIdifTMRegpWySkF/AU1D9n6duWMh57E9GLm/Sn2
ckllDQxklEojffFDd9m4mxBqVXi6zSZ21WcfBoVesBG35Myvj/59cN9m3K7JkK8bGP8UfG0CKAyt
vmd49meCqYrNqSvsXxkA5+YLw4pZ9075iLkhlMS8ONtGgq7YWHmcsUvVdFbQu7X73SHnQApL0n3k
SFjTLeukQZywqm7CFhvgeE+hNzGz/YZhSjkwkh/fbrncvmegDhKoW+jqTnKwjK+tRUR0kYloXb5y
JDkuAsmoDotjKGgUg0US15XM6C+lfRSaRcD31qUd7EnkYqJ/p8DKXw6BdddgIRk26T/9UImbztZ2
2M2HGs7+ycGVJ+6aY2MuRyoFBluzi0sk5hiHl48rdcGCVHzYM42is375+OemX+4qxoC83lSFh2IU
kQuofKZoF8cGiHCzezC2/MPMGzafgitzcn34IBnWJVpAWkguHnvkmhFKsGQjjoANhdB/mBL/QBJU
nclw1o1/6IHgAKgW0m8vCY1knKaz5fkUp3/P+JxZbZUOT9q5oVO0jFvpwoSlwMq7vnQnnPH/DWCQ
oE+onKuiUbMOzh4k5i9ByyoYVnqNOq4VOUSgpvWXgEqxvIQZy0i5BTNr8kPMm3GC5471FpePD3gM
BUG/qUBXY4J4HWTkV8K2aF+8A2kfdhtKs4dTzAOWq9B/Z8Y4t0npdr+vl2tFZfI/gheBfBXP/mFU
EO3mhWhTVWHMzp24yXwmWgHH/YqlzKQKBoIN3+t2A0Xjpg8jmpZWm2HTUHjwhUhnQLWDdBB2fYYX
CnV722IF8MIFzXI4wYzpFj2LkSM5/ppuDGneAKO19J3JwoCHopWv1IADlFIKw8SZ+wxGUZxMxCTS
xV1u/oWaOGfbQauB8lvEUCF3imZfwSiyNBMVLS9Q7DbMGwDTTHCmccnkrCu54FLBEZCVnEWZNrOO
Lros+Cok/9grptGipUTmTG4QW7/OMqbwAiL0IRvzAzCl5Z7wKsHEMf0JHkm2P/yUDzTQgBqRZF6n
7Mr3GJ5XKtKb7WT7XU/o3NoQKH/pFH472pY+SdgbJ3BgJSC7XIxMDUw4x00wRlxRm4J7aXmIEqKV
lwcXPwa9uPQJG09GVoqk1WyVrFyyvN7WmsXUfPXf0FM+1xO9NT4/yiy3KekozeDI0V7dW9t2ES3l
JRieIdc+x7LaLt/S7RMsDMzxYZNCwGDvhdeoB9YBEspQu2etm+fK5f7N/Cl5v6hV9IC62qQzVKT9
voy0O+k43rVKGl4vQQCzxOAk3KdZf2i/d79UlM38J5XDDIFa4XJRVqe41nquN2r8YnFTK3WcnrJq
QhpW7OqUj+qh1c97HMpibGfPtNev17GPQcqNm23ZbCW+TezAG7Sg9sMQSyUXd1KBIjbGryXrbYTr
e4xEsgW1bloh6Qqsjn44fsD0yRpNItlRYZrB5OxYt3zjO77axQqbi2C7IJME/R+HbOqyBEeDF1xJ
Ywp+0Y50KcR7hCDT8dfGeTG0pk5qLOak16yuLHJvoW/bFu2LCDixbg+Cuka1sQbHMUH/z7Tk3X7u
vpo6xmola4XyA9zu0ZMEmUj6I2qU1HZGyoPa47wDpSyixEC4idZTRPZpMlKtZor/Hqm+Xxz/wvAT
sNSpm/ILsH4Sjko81JA3VxfWWBTqNvYcnFLuKjHXc8hJwkoCKCDC3FRRAY0mBmKQFgZFlnANpybL
6/CeHZ+APL1cU0HvHKx5sKNVIN+XhaxQIJBxZydoCcylgwJzrP3jfWiCZ++byjIIa4FWJpD7cQFP
V5yQIq4T3iEApE+LM8L97i1qsi9aXRhFK3Ynl/HmR3lvct0tIzoVdFUBDyjvURF4ThtZJA0+DLDc
b8K2uR2VbWkzs2Xff28vPGV8W+VWl7uYhzFfZwsS0PwWViU7L5A1JYsmO3U4ukEbw+V/1fMh3oPl
d6N0wyJ0W1gKVm75KeniPC4J6d5tkSe8e82r3zRZ82Xs5eGGP4bE9eEtcSJv9EPI/hSyzUi6RLmq
VKWSHG+FtlG4juZLylr5siMJe5ECpZzcE7KqVASRSbvLevoFIt7UYnjHeZJFOwJidlVhHCxdStm+
NLaeq+P3XZFNp71DHgs1K8DID0gTLx873rMD1QU5Be+iHnVPW8DlEa9EsT+1Nh9r9Lx4VTTECUAp
T28lwN4+Ni0do3lW4KsEFc3+grsnhgUK5/TDx0oczAv3ffOoM0T1C6jhxQQ3bO+XQxjMCmyaswhe
pKAdDrHuacpzmFkNaS8rT3UOMoiAE4DRNtxpJh+FGmob0wTsX2VuZWvzbqxW9oXBA4eCdrHI9coS
dQCzasX1VWsgC1Ut8YBM1o8LP7/byrKlytTvxuGogUTOVq3UNJBElOhDiahvkrjqmidY0gy3lAvg
IxJyty6495+JcQGTEYt2c8aUsQXpxkhBT4QdoB5aAhvG0MYUoFuIECvE35n7nuactPI/uDesaGfr
BIVZfPAKxSff/TVTgTHcgRMFEjxzTalA1sO1ZRywDm8jchm6QMi9i5JDKvKdJHKL240ZPlBC0n1o
l7TxgE6eait4iwa0Zt8ACqD3m4PiK6HOJY4KgQtC69Wz9f5Op2tTwgLRbXXqLcIGeMXZS8FpIdq9
K+aB4dkR6j6vdxRFjQ4RVH/rUmDZdaKY2q0Cj3ZYf+IPa5YV++86XneqNli2K+sGa2/SnvbqFJdP
CjfOqZRI8pC2ifO74pbGW4rkQyl4tdlpPe1JHMTvQTaBhEi0oXTPgI2Ixn5SbdlvF4nHPAUYgUQc
flI0vd/irpNjs2DGYLBCPmLIUQ4gIX7RPgctqThRbU9j/OnchvSaev+5DY3UQK5MqK+zURe+uuJq
YGDv7IGCsDHIGbtTfj9EkZFmm7j7VRsrJnBzOtLvakjvJYxJBnhD0DA68wQ+2wwDf4uciLGGqzTP
kg78R5k5RZctfiyZt7ejWqSMJVFEYuSSVMRb3CzSlIRFvRzxGQVXDSmswodcCJzZW0BfMRPK5297
+rDU5hdY2u0pV/ADvKHdeqhgqsPqfkbCWZsgg1pVdWSpZ+/tPvo7gaAZssGhh403z3JkPzEwf+ym
XRP1gXsQCCJ+kZypkuaPfG2Epq4dLx4BzgIW765X9Zb6T2ugJQIq0Uyj5Bky3wvlTNcAYhLX/QhA
PFp1Ea4GS6Y8tHLMfHFUhUR0l154twtK/9KK6rZyWRtvH0/PLjBJXN7Hy3nt0VDOJPY4F1GBdWmG
5aOGTAy8zQt7bWt4m0VlO7xBsdgSI1yIS8nsyclPzUpUzgM8SvKI7q6GMZPTWHjzhOVRjBymddl0
2sXFcKY646ybCzL8EDqp+UyDIDcB9Q8G0iMptanLlqyzgCd085HAZ0NIEgZoUYjw13tsdMT2n9Tv
upkPTEb/BGEmgOvcgS3+YtG6hQpmj4nyC3VKsca1TQj+wOJYf8toXKOfxIrx9d1VUx5lxUOKnmWV
3YR+0IgrLIupL3sRyICdku8mC33dnm01SvuZFY8ZnraGgwsgNegN+jsSwHqtlMrOTpsU7MssljjZ
Ek9TklTL2N2zQbENmwLES4U79QfEXRhifpFSbB5gzRNfk/TyPtIQeS5WOybqYU+VJr2S/bu1d5Ra
wM7YzDpN9CX+y4kIuU+X+U0b1nJaIQw0jZUNBL62oZSBkGwEcki9NGTg43i0BrGBcsxphI4qk28a
faiBWqtcwj8GR85qoGFxTAE0BBPhGgtkMpr+6Gea4AKcUAnkpysVrprScfRpH2ot8GkkvdTuj4ve
3aDCWHkc8J47LGZZm937M8ZtSj3XtHmYU4JHlS1cf4hTGo7lCMNyovsoqJ2PCK8VOUcms9gh7jtX
64w2CIMXL3rWohSFvcwdNR8JMDYmfcZMsuOteEpA2IuLSH5kx+7b3xUc/o1xbT3/RaXWTSE1+1DA
z+/eqDf0sEBu+AnReNSlB/OcQLJgYdlPwtYV6z28SAJoQsFVQEm8GXahc0N5HKS00R/LNX5gCiLZ
gq+TTS+3vsgwR7igjr7J0QsNdaZO2UP5j5JjUly4dPCy3vk/672l42bvaw1g+drFTKugi7SYg4qn
C5V/D9ArkkB4AY68Z6VYWIHPbpAkS/xudVv1x+lDEGB6OM/tn9mLJYi3PeS77EfNsYyUxj7Ybp5U
O2K6H/JcQJ+ZswygODpWKl6OxJ3km4nkAqKx/2dCkiRE334wBism9Fr0cMTUo66MKVne7YUHB3Uo
54LYiIxvpkbcwMu3LDEeMrNtcd4+79RGD4xrgCGPQKKyHuooVGZODOkkw4A1zIcAQD7oCYTwC5qI
8g/C7PCwDHl7vk6+quJL+Vi4GRkmNzuyfRP29LhGrVeoZTrMfqB/y5HuntS7M5zuDqzsJVteohJH
12HRQjR+4HwRyRz3TqZ+8GIjF87gpH46H0rOSM332a5qrwPpSEybjtaPsroZ7nnVzTEBdSazVzYZ
XeboxE0HUIGTUYryfludgya/+BHkniPLHQqciu1vijzG0dmPerU2Bo8MqCKXSfQtOJckkO0V8HjN
w4RTESS5sqHPikrbqakekrI1IB+ZQy4DFRuDl9ffNM3AllIY9QYMJxxsteCY5CWinVZNbbSuPCSZ
6Wg9Fid5eNqom/IgwOaYvT1TWMkuLlTtKzCEm4f4FJmmecXdd5yC0UxuiwvIBYPIAbLElVfcpzx1
ABNBfrk6ToUP2bIMQWKXqrd5cN3sZSyF1vCD2m6gZiccruxbmMJ1+juz1FALMqrMiHD0T7N7UXMC
WfKdQbG/gMmYKFiN5Vn9fGDECk7gw9RMtMYc8O12ZUSZWZlhceezhasgWTicf+QDD9gxDZoeYSgc
DVrSNJlhpNhudRQ8Jgz16bBRApr/NIWNQ6ceVZWB1ryA9oFUw4WK0NkZhdUWvslOSxo1h5QuHWo/
U+STzSc1aZL0fvdsLDEafNuUjlsdHFwsrPOUehlaMvIOfSfA0ql3vjAMErlPm1hebIqEnBfwsJGm
doi0lZK84aYj042yIRz3W0SRbFd3ESazwg0FY2ZZOi9d6IEjHfuqnAtXDL9fF7JWMyYipwFmKEQY
L2ynRpf+czCSp9aPzzYUlJYfo+XpT6BeD8uUQynE0eHHPde382nxVmpurRu11eGKOdB/r/S5xdRJ
z7VPeMIiq8EGo74pYoaSRpk/ZbklLlYqoSX4UgnDe3xroOY68S6CRmbXG3I3PQWsK6UI4UfI2kx6
IGjy3eO7EnMIQvmeQvbQolHWECuNrXt4gYVdlHOfObbNr9874ibgIS+9pk3rRK7uc4hRnr06D1+k
WIoXHb+GUPVqj23DjW2/EJbwXkE8cE+e7TBJgVoAcwDOXRiDrk0irukU4TDB6tYI8jSe4JF/Pu2b
2APeedGn5jaK9mBPMuwC45w38jHl6+JSdvo9SAyAgRFAKOtrVCywK5h2zzfR6mqk84s4bgnyuV/M
0tjnhJljuySQwPXW5W1qxSmDFmQHg5pYLAGzOnGOZJpwDo4T4V4qAfbFH9UlppxC7i2FDbcnGmO0
Lnpnmz8z2mwsqY5XkBWcdg63Wxa573whCfErYgNiOzecuheXQI2KstozfqSq/9M2qEcDDBoxsnwU
t5DLykMdyTOxZLlIegUeWra1QIzQVpB3nrHPl168tmjAyXg4dsacxvv324SUtCp85XKevvvI52wE
g/g5dLbQb09GnSzp046tBNpOeEkxH/gjXIrfg5w9X0payJSvDljEP/saUFIZP8aHvtUzgNmpZlCl
JX2U6GAj+hMFzniw4aPjFcEkCuKC/Fhdy6MWNjVo3l3G9jkYsfgWd+/Ttm8jYNbJ3dGp2Pwlwuo4
M5kzz0TJloT0Icg/6Mm9qCRs5HORnRR0JhXbydVKWW11twyeG7cJU0NsCRv3ZSP4Yaod816aEjzZ
MvebYIal5BmpOyoHsZfVBMTEPiP6AmmicGPB8P6w2XTRXvJ6anymgMmabc+RNDKL2prne5Lyops6
/7K6XrvvHGq4TELPBGksnxSbMjS/Gg50V/saEbpUtfMwS4KnAz+ueg1x0m9Un84LundghcCHGdgJ
0m/2wp2dDFRfztgyTlJ4An/WEgo7zGqM7iUXL3R6Zlm1QWQU4Zipb8PQTFm+rl3ix0uOonnXqcKK
manNtgdfUlsTPiSp5zH4a4mzaWg5hOoZwe9pQqCVWsZpM3nrNVCRPHXq+8De3ErULReEdpFpHArb
EA3N/5dxLkzRRODGpNzaqlFTVhbzrtR/CWf8p7T6ZcTD8ls0/uanYTv4DoP65YH5C6xnEPaguYL8
25qENXx5/FTmYcudb/vgGcqaiR6Cn+s4m4OgV7NP1V4ayAKgvKlU0MHPUePe7odX12bFoD9cdfD0
hz2oDwABVpg5KLw/OBcnQ/J7k3QQKiDcS/iLpUilqU3CGasNRDXDMx1KL2Zz6//oa+4okiS2qK4M
YDy5si9xsAY7XNKh79yz3vEgX9iZK06NH1rD2Tfv3fuQNS+XCeiF0WZY2pVSEBKfl4gTXOwJmOl8
z8tyvBdSkztng8wIRBfBPTZvQIDnwc6Hq1grYscL6si3aeXe6l3k2K3s4yhWCFaQKR5JQDcvzzuP
YzaT33StCUqwVc69GA/Aro2BGlOYQAS17XmzW6s492DSB3msFD17EIno0PowaViya45HPxwVTl+D
8CQxVai4zRqBf83SFgD1Rk+vMFbrhllahKKgkfY+6IXBJDrHKMxiPy1r5VaBjq7YiEL97x5VxSj+
MmQXfKcFVcVLtWhpIDmQ0tj7QtfczPIXi0bgqcLe0TbnCOjTlp+xLkPM379rvor5LcRH4Dr50k9s
cfmA+XSBlee28xXmzT6YcsuFr8vRStKwXlvXYrMbb3anSZSUuVIDMkf2IaxrxgOCuRClE3vHGis0
O2dtYPI7DArXX3ul42J+jenInUKEjVq9s7mKJhT1B9+0LcSxmNytll2utUQ7M+kIe7aaEzXhwg4j
45b2sGqV3KPebm/ZtFle1zWOuUKLSmv7R4QcQFV50ksFLdAr6WAIMjBndldU5RmFXbWvWhupXngN
XUoWSuKJdoiC10HPbQVWnrmXizTfv3fgTLXXgtKKBjgCnkktxYCUpcd59qHiYXnRWijiVoY084dP
uOqJqfhpEkATCG5GCi2izNO3kpEBwauNcM4Gz8zxV24s/kGJFUVxp25HVeoqI0/+skIsi2ZJ4mG3
cbnLSELaod4CX6CHnmakH+MLvP9VPlDIP86ucG4N9aMvxfWeTxTMydOtTiZAURfqDty0bYSZL7RC
wIIthKevtVRjHHrsOlETxF5+gygg7rQ+Bc5ArjJRWXmnT6hVAg2brr8aXrGsW4Apy6HRcTxnNJkT
pHR2a1+9GztTuj1T8XftEqmGxuV7oTQ4uYx5Ya5W7QsR3kNdthUK0SbT9idy8l+KZcBv4y6Tm3OW
OnggUG3FhXkfz6ITt73N60Abbfj3CF5nJi4NzAsQwMM1h4rOEyei+52FWhhTQmzUCgzqWJEiQFp5
2dLzVcZb/pMok+87zMNpCtb75lrLUv192HIzM38fXeprSjTfmoMhfkAfi0p/QsJ8ylVtKy8Vlpaz
o+D6/2cD4/0E4EbaLVpuytmKT4MCV6KomdsEvB6yxxSCHdN8Qz0q+QR7eWKs6tKelHAqdqQs3QAg
Ix1QPeVYvX/4H68PiLPIMrDDmwF0NlB70X7NGrvh8LYP93ublvXJYzNcAxaxveAbfTgsKE9ofk/I
3Y0dmRM0S9UoFlawFIO+1KjJL40OHbPf375NG9N9cg5XV09oH/oq7nMpNMt7VjSKwOHA9KO7qd6N
vd9FuEVxjFbND7hByys39hNkkE+CstAMx6iJITycunnUPfxAKg5y4jJqxLoxG7M0PBUL5qLaa7nh
lkeDbxhMn27cpD4TW74K7Na4YagqDlzwDVCKURsALJ6ijTDLIVxA61kWCCknYT07m2tbdH6uQDoW
EolvTKjGccPG43MdzjQfpHjem8zCUWG6KeFEeXgvvOOxbpPHCvzOXaLM+01UfTXZNN9CjWg7LDpt
kbaYRJTu4yWVpql20TzmYwrNPGQ0DkW7sxgJ7W53fvsQTCkOe75qS6E6HciOfFoQEmp15pgngRcp
E9lhszmzCZPw/vBrrwEfGlbzcbvWFBQXbI9loNJsutjbWwQdLWnI7VQ6lzms+dFNNkcl7Gpbg2Ks
ftrTjmV7onI6BLy6OnDh0akIkO/Zf4DI5ObyWb3C3dPH37egzULj04BuxJEJERXt3y5HnObc8O90
owQ2u827SJhKhiE2S2jTuoNuhNbiUdwY4W2yO+tJN/82B6E5JS9JK+14bc9ZKrFp7MPhLJY4h1nT
7g/cVu1WJkU/QfSpG95q7ERFGUvGpX2pqLAQ/aoZaY13C7dPFOzcKO6vsqiq8yI7L1Ubhn7/DDNt
fl2LaT756q0sqShT10rV9sZ4obczjUNTRI3NjF4bY2BG+tbhpqmlsnP6K2/t7RaE8jI0xEkL8YFH
9ePPeg504rApRk2DagidKINI79soL9Bb6fRi37V34lSwHOp31wtrTs6Nx2A74Z5+17otK0FSJ3lT
HeONOuDEeW8sJpR1Bz057zu617p3Yit+YzuJa4fa2BVLcD0wsBlE71bgVtwIckit/86XmW9qlnOx
U0I84HV0vspnPgjF4Nu7c14IQgNK28CI/0QVPInkb8yXtsjhfihjyF89TwZFY+PSBRHd6C4tpulm
HRSbOdFTecaikTxhFR/Q36I5rb2sOo24kYrkEz6y6AJpYTMdbxUHVT+hzBok0FzeUGj8Mr/SZqMf
1zhlEiC12O1kvJ0kzr+17x4myMw5AsJDEtW3twvP7+5k6dcEx/NwUN57eIsw/knUA6sexUMB1SAf
BWZoE7rg7KBPFvILJIZGXS6iocGFal8EE182M++4ANo/YLt9QMzcofuVfjXptye0IIbGyuFRC1Gb
bIyWYEmi0lRV6jSTULhg2z3imfnNDbmTrN25gJgZcmZSW+BYwIaxfuY24fE9oHLcQWKXnlUOAduv
cTDv4HpkSMVGBZv1h9E73iv7isK/CvxoFYBIYOe7fk7m3iZDGJeH1BQqHPPj7XY7/tyNiZ9K5PGh
z46znvtixJU1vKNdz6CwMbQa36gnieEbaC/H71Jvc54LpxP4CkKqjpG6+a468adJjwEEJ2XoKscC
pqNVn0pYL40AiyA00lEmd4Z3ZbbdsYpxKiDWvDgJjvkebj/EczEhbYx0/H6dtTRlY1kgduWTy2h4
igbzF5sISTZkKzHghtm4Lu8NXH3n1+rgoRuDAzw1Ho4KX1SYcl3ccRNrz0luhlHNbW+ZBG5oaCAg
4ECA1cwUFi0EqkYpWni26fOhVs2ORWsH0Z6nn+XDsZ8LJVlcgEND3RmGdhfE9Mjcjg8zJQsV5+8P
fheqAgya218foJcUqXoZ5oB9xWBZorKk1eEwRt5fSkYrpA0rOC19TypLl0+1wjpjnDOJ3auN51YV
SyPpaISeP1LYrNwUZ6apd6dSG2RtZmBPr++6z4TAm8muF4Wt+s4mfPZl1cVbHwl8eKCkQ3iHpBMR
bM6FHWhAfqvfx0xce9E80RSa68tRPZWwBK1hOt4f4lORR/M+iowSw0g26b1UmA34AsnzA22GHoc6
mwzOe0g097cQJVxSO/BCaRHxC/cFC/AnVnh/6aUhbBZv7frJ8f6TLODxhDFN2Sn94uPGPM5R9Cvx
ug0+fTvN1duB993Nu4Dk9CkD4ocWpFPUApJCFKkz4Ng5ulVP3Gz/eilwRbVrVPVRNudb95mVBsK4
9asJwARHq1RnOFl2YPH37Ct0ekT6+gF5t7YCtvbKT7jRt76vFkg7kySgWCkurqjCzVAvMJGAzzyB
HRvJfVMCBldQ+F+dAIfCSOhxDvchm59eQ7nK3Pk784eG30xOkb+Krs5h3fEhlW3oTv/qUMrzOumA
is8MNFDlxxtjwggdRmmV8lSQUvO5HTEcUn8CTbKBZvelKTTOyBOo2ybbPpNkoYkVLz1xe7jgdME8
YHNBkKz2NoyzzRKSJ5PzW10x7FK+9GTKZyRKEu5pgJ2N8hknimbkmUreRuFvXOWhlI2XNs5EQytO
sORfg/XoE12gCOwQuQWG/G0gsvp+5fXPegnLoF5sYmYt7tfwWXtMeWYhIPlyCnh58V0Drxpyhy59
PEqNFKiX1QvavMeROAkHkJ0oY9TEiIjl7wNUT7vYlzDi3XVyRupNpdzM46fFgpm1VIwre0GHBqVr
UuaFpZGYsDBxLL0j6SAEz8Y11ug4FeBWdfu/NTsTIZoDJAwFlN2ViuiwFBiqPVT0HSjgK4a0gqEU
Q7oDiE+x8k7BDUWq1DE6VJhQkoo+zC0sQ+82HxfDnPvEpsijA4NTPAeAjewQJVGJkmIpyLIO0JDO
YEi6NTwUcbjcL/BuQYlquTB1kMTNsT39SqMmUMHJGhrZoW1CjsG3rb9EK/iPvkjWXmHLbpcKYZ7o
Vt28Hh9kczpFdAmVteN1ny5Zpoy0QZm5SOVYb88o1eD9zEmbxR0QPtZii1RqqihK1I0S+uLP8do1
Er+UV+CLgY3n0YaSkkP5iLi9qvolirr/qXVocUIdf62/1quzbXDV5/PHNmA2Q5M5qGapC+lVg9e1
lqTV8GiEl5xYHZhaeO/fVaT9PIP+vq/OMakp2BEwcTTE+GhR0+WppSCsuHLQXcMVHBha7BoYTHC8
GrPRCQZOwWdCiJKdQ0tD3pBRD8Vf+sh5g34xwTgCl/lhoA4Y3OdXV8xVxMCo8cxT4IyKLZju6cgL
VXh8r3T0mw9Pp8L8mg942QcccIjeBzWbLwutNjRIcFuhEaKOKIjy5X7xIW9lZow+VNxdLA5fcsqP
MUAe/NZmJGPpmAM+718NI4eXMyd973R3accz79SD0zqKjiC7SZ6jqcOlVG9J6j8SJIjQpI62rCVk
gzv7nJ1nY1WKh5/kKHhZBuwLhJviOrdDbNQn82WoYj9VXPWFaPG8hqxRbDhsgMs70r0K2trRaiaO
u+AreCUfw64pyJeJkWV4J/R5e86nEh/N+yBJ6Kzu0UboBMz7kYxP7/b5B2cL8PSeJnUMR4/e/c3O
e3Qf6cGgMpvgrQ5QYT1OrOatmqWAYHLlsEteC/9518ylJBaWdxsbks5dI0WQdBdDgpkyvj0Kug8u
ok/4Aj+zo7Z3msoZk8y+57HOT35/CabS8fvI5m4vJ8m7dMi/aEZ/Nrg8CWZUWp/TTRASlcGIyxiY
dDVFK7FBscp5zUTU6hadg+HBtSUMSLgzAusMzYPR+bdGxXueqmgme2LewRdXjxQ7PppNYWmmCAZf
cwMALTV0su7VSacKqZ4YaRLUNpbJ9Y0t44tw8khNa/whDiiRI2UVNkyE6ND/Eoj4KZIjU1sIubN4
tqAx3r5kdl1BHVlYzf6/Sb9jjY3UQxA9VYKrbxoL+/7XCi/TUsMh9XGX8e3GVI9LHFy11q5WBisG
9QQSuCjhsm5hhvnrVG1ehzrp363uFzE87h+KwjlWQaFoR+zUwhwFoZb4xb1IRxD7s7uaarAzBA1x
93QRsj1y3wUEy4nd6BlybUnJ3YCCDvahULAiPpIu+RPMpl6lrdjvRCi96D5Xe01JjrtludDBnGii
dAm4pMXxaLEBtvxvHAWvF2fYCB+MzS3grv1+guyyU7/6LapeqnTVUr2BE4EJAysbN2d6Xp5c3aUN
GYnk0jqkmALVAMzH+TAnllx881I22Jb2msqlPlFkQGS6B4EkmT3vJspEUiNgAgN5oSfvU5zshmPf
pHIZzXnH08wB5WUG0RPoplsoZXTL1dc/huiDThDiW3udmA1Hxwz4eUEFuseKAiU1xm/SBFZYgx36
q6Cs+YsVnR7otX07G7rMhSYDY85G3bZoLmgz2O26ZCTY3ZUEJ0wcK+zsMd+x+JhJNRmFzT6z6m6R
dyNfVdJaGP2/GmHywnQ3YxE90Dup/TkpN2h9dAfFGzdcq5wIFNPoIkBDGHENo9EatLxg3sHdf5tV
zfiBcOMFtrJ+pGLBwgUBk4wQj/JnYrYr7VqA8oTcx0q6xr6Efoh7lWuakW1hikG+qn3Gte4mnrB3
Cy6padWuUIfvW08STtM+aO2AOtDta1ROod/CLd8TsGPuxNuYl9ihF9hkQyMnhtxP2UH712bQ92Yj
8Pw5I36hCHWezn/jkJzo6AAH3j5NRkRbugDJSLCszXUehwiwcBE1AFEdRVIfqss/EpAteUIw1kmO
LZNyhHAXbfiSzxq33SeCJG0Br5luIek8e+OXBeah+XEL9+mO7TbFyjoTuYRrr3xODTNfRJ1yXf93
jsTXcvo/HgD4PcaEiFf2UlKvJMy3UW5rI5Ufx/7q1LEDKsIySEmYlvv6xAHMaJNxweJrAbGRSak2
eN91/XP3SGxEF0GuFhm+KeyOa1XJ9ZfEav2JFmTsMkNTprvIdhwAXmCnf72MtojBFiwNey8+gS+L
7hmZMS9BpibU0a9RIozysww1ebKq697MyxltswdbcANYa+Jr/D8TjptC6Fc0JkOPBSZUdUUKh/kZ
9ADnHHo79IoapyhjVIxU8M2MM795rJFBeO0M7z5qm05hiP6iWHOqw9gTGT9mcwSA9NgBalhAlnfz
WYXEO8dE8eXJ70mKtF9F5BRlXT7kutWbdb1AK402FC8+u6mwOtazDFpCKcS6t7WSl5HxqCxwj5Jz
iWG/Gq0aVLNAJ/qTqZdV8BN115LHPBCVVxA0m0lJ8nVfj9KTCxj0lCqEWn2gxnn3AordM6trRshg
5O+F81erfAm3GQf8JN0FgoPElA9NLkKvRywsT8HruI0AUvNnRvEXWqTa72RQ/Me8+mnM+U+Paqq5
Mi5LpwlByExwfsBE71qTiFI2Hd4Xnf7qx/IKNknwF2dH+YYbIHA+acs8OvvQ4qGiRDerscdcX1Am
rPZS1OSQ8KbGqF0kABmyyNR7Z5GXDKnTDjGiqtG3Thh7CsATCAG+zr/HR5UuyAgfAtm5IPvlrqRT
EdNs5n75Vyu+iYwAJeCziR9fxtKZzEoC9IRQ55bCIASX83Na5fe057rdvsrcSzj6Mn7uwz+hytlN
dzlbSI0Q7Eopi0l3lZh8I0QlA5Bg0VC2TiKmd0jdZbdapRo+2xPFhLHvebVXUz77aJ+cTTbyL8d1
tU+90SUWdQsxJiM9CxM+vhoXyr2dPAInpp6uPxGpoYWKbx5r4959GdnP5n2tUBArspX9Zve4/n70
DcR7m9StAQeLFbfaS2GaTroxTZz5q1KfaopPrafR33RfVvap27E6FMV+dHNYsaA0zhQVhFKmw7nz
sW7yseQKtqDRu1AXyBidZsv6r8I6D/RaBquUb2bclGM9I/Tywm78CngtRgtXP136cdmReoDOtXvZ
xGkKoNmfCcFI1Vv6jP57n9t32ZR58xSKIiiz0JpZ1kBFlkWNt0jHtVqWYvf1oKu46uVqCEa1HqCm
BhBFRT/zi9NBjN28UHvWBY50ZRL6tM6zk2BzoVyZqj7iJBcoWgSxDqMHbCEcfbJZOG9hrzUEtAxj
HDbDZjO3bpRDM+pLqmU1jaAWR+IxZ25JD8UMHxxBAxQIeyeTrthJmAydlSj0mAVmDXNsGbun0tO6
R6nTrntiYgaEMp0AeuCMQHqvSnnGRFTTDPGO4yXmPR5s7LH7n4QCeCy/f3vXbtd9s9zPskshYms5
QkESjSGPDEdJtuUu3ba4vNc6Uv/nVw7K2nXBRoJK0iqR0k7flKzVyn7UfPcyXAOIOPg/vDtnPEtM
TE+a1ncSlc/8FrHbEwsHY2NAjfR54xP88hAJ7yJGFOvutRYu4GTdOQxAXNZVHvsdskGCFj8Ep1iD
KBEKhHAHxWxTlXijpypYcSFHOxXE1+oOh0xFP8BwVev8NLuyHngAcCU+L/D+d+jm3AZe4BouA8iT
Pa6UOI7Cu+G1y2bMkbrq10sMfkLrClj3fqrkkreWWPBmvsIE02SAHRCeGihT3JBOTsdlSKuMxXKH
Hzmy1++jQVMJiks4KTVlNjPSIP/GGjcagcW+Yua9af0zKd4x3bnnSDI+3urlajENLt2d38dNG3Jj
PFsdGZcJ8LY0+1/wnekNly0g7zGUSyIlLc7VIgJ1+Ew4hZ5751ls9c7odQGcPR2RBf7wgP7WrDZe
EdVVbqskr85EKVD3fDY89htkNyjNpcQtxhCUU25xF741tVZ8y5aWub2x0inyOr6PPjMMwNomtcdJ
Ba2FP/5feNWA2LASzqbagwDH6CzxhC8CACoUcFkw37p1M0BtwnsnC4lshzoIwuh2VYKovy1bMa8E
uomeM9BLeIpN5+wkkgPVzxtmm2pMZU6qSqXEgl9yO+UJ2Zjces6cuKT4sRgA7Kbu+Fzs6JdWF50w
GRpPBlj88AXFPGERRdz5dTQRym66IcBUgDJoeyfgy6dHSR2/V/bfirqvdgVd33xuzl1BMAHhSmdg
vMxC7Nxy4tn+kywra1UQe5acU8YlWJWGOa4AebugjlTakky9Wc7mYVC/ujjGoMJ3hu6yRBnUYchU
5LUoIoon8CZ4mEGyYNfVNJpu9y24k3SJ1ghGV4BVWPYL+MJluqOi+jFEMyijUwoHqaRRvsJnrr57
dzo3Nu9HON9UfwzsHO94ngOqypoZqDeZQbbUorP161NG8n3pr1cWwYhpbn6yhZTDTD2CBd202RYE
bpyZ1LlKF9cz7+D916j3E8hZSSL0xmM7luEAaG0xFgjSFnKxKnRO2FijZ2Bxx4ny7sA15/WNOyU4
2xGixGkFKdVPaJIOoqbd74DPUL+IooWnkmvWoZpj5gPovg0NuZMaRNRCmp9cZP4aQZMdAq2++DJy
rZYKlodTVaK7nrTcjODN167IIZjZ8a6YBuc196eDs1k81THcPenWjmOkC/M6e76jhk+ltHfOzpdP
rXjeaxrrso2CSdW5Ahgqe4NwpeROgyQU1dlavFsX8oo4R0TEmQRIKGDfVrnPjvh83pYwL6BuBpSl
pDeS+oEj6PEBhUnx7SKQAiuI97lidkmcbKFkN/n1kfV74ZtA8UXxCkRsKOjmz006sHBgfOJyBqu6
/3Kh/52xXAYlAwhCDbTV+H+SvYcBYLyl4e9g0Wx6yRGVQSPXSiSABg9pDmiQyEPJBV8Z8kkd4sPb
iXkYmb1v4o/LwRr/6af9mukQgVz2XsHVeVaq/sQY1m0NnUC4Uz80ZNlUfwEkAnwdFkJg2A9o5z56
o6mwZ4ROvJp/XHKqN/7Yii+6RukTc2OcYtJYQeSKstA31V7dIC28Jgm8jqSNjdosbBIhDaMlFUvd
7QCcpOdPSjX3VgTG4Atq/wYmdrv5w9SbROiUPRedUkRsKt8tuw1VZI8tOiy/jdx0yWSmiIKF4hRv
skA/aKMA6RtWSEgelZBsJXKX51YIHM7MptETwaaD8jOSmCiVX8vfTXWjx/N9oao1BftRYlcorBS0
bibEX2ezyKg9X32koOTQbP+d/2Dr6YLVZclqQjVa5jy/P6WXXh7wiFFOefBXntNmd5KjOzPYB32h
ekmkL+WMqpd/fDNLus4zSoQaxxUfcJduAI0nXhiRkiDkhxwV2dpgcqybvA21rBnVpzRm/CdUcA4d
+glnXUeibiQj9ExsxV5C0BfdKsC/dfUm7EuAGM3MJ8l8F4/a6r5SzojJ0H5WriWck//k4149ZTH0
liZ8LdvblIOaPXvBnj43JRAPJp4ukrqBMDtuuLEgqSvF0R67MbMzuPZ5QiY81gp+LNpdUTvHvz6q
o2JZv5WOdjMef53EG+k2UX2ptIHYPJMCRQpo0obTwxFyxzMkpO9QQsNvJidWo6MJjpeLvtG65sEl
KZBfzQu90ZAddJ5CoqNNu7peEbaInRWfzmvFId3MA2w6tdFwk+f6dbczsgz/QLDEvs8CFainMbfs
bYrh9/7lWyzk3nnREGtyhxrXtslBENsb4UX2buq0dEIoOhZE9+DvzZztN8T8MRcAKhKt7T9iuzRP
DOm0Gek84O7Y03it2j88PfKztko/71d5GE4NYGRDIctf4HKIIvsUL2jrcOnOwxXZb+gp1TFOAd7x
MIgBQXUs/JNYL/gRhLID/kAKfEQdogeDNIer+MKXtV6JuCk9jQ0++WPTi4NWJ4kZpGg2invVebIQ
iAhLD3KiJDSY/H96RjkRMqKYsEYVZQsoT82cZokNsLcYQ+iErm9fc0aeZkkp29ifhoIaO1MIMbDw
ypdqaKagI7Ni4bhotImNrjocQ/DwP9qly0dsoy0eEQIy5jK1302UyVXfVwNO9qboCNfpG/LgQq3Q
9FUQXjSbNt6FWWHyf8nLSHaxhGG/nVYMFJ35BldVvoxqu9JoTDrDpVjmqoACiBWZQYtgBungp+ih
W9yliib/K7kh9bdcwAjeYwapIprCqvDJxeieOWlbfiAOs4ovlQZas/ZtPZJFgDoOPlZGG1oUsDwC
a9Ma6VmKFaY13W6AwrQASyE7nm5ApY36sXeM8kzdcoxN6y/u0WbkKV4sQhU2MsDjYmzR7bGT0KH1
dLAD759sZn/DKn0bUKR29CoJ+r8O29R+RbjOwnYnWUhlPQz5tmJMNWt6kCjyeapf74uS+GvaQhX6
8SgFIrAjGEu9Lb60xelan37I7wQe079o4oRpUpW1CbFUrP+GaIFCgIqlD3JFt6Ne2i6FvZD4KVHM
b3rSwM1psTYHePBNn0MoTdHLhjNpkACTMfT+qdfOTc4tulIo2+Swlju4IVvq4tNewtqhesEQBFM+
FZ/5ZhaYw9ddhfUgwCZYdrLjcA+Qv2vJOsoBpVFNG8FHeKHF/vq/0I10NbX5CUQKTGG+bTIBFHZw
FqmMra4K0P/naH9tp4J9RztQ1LzkuIdLTksv33bVuf9eNFn2IhjBAoEXIAOZ5ezBaZ83sbJIjD/G
fVw/kcUxl5bxiO638FPHZ0RhznX/tuFItLxiEnwW2xcFJ16CUPdnoqbBKQoJ2gIiLKnMG/0zxI1j
fuXZPKQioZRTzQbraTJ9xquehUR8Q6AXUjvsGD0CSd6fE6ByixtZEbxQTkb2pVYZ4PsRc2joEI3/
ctXHQxXN8D/XDqJ4+NJx/6pv5ws6V+jjopYKIHvsJvy21Z2sEpD5HK9BVkX0aHgNFJ27LcTdCiqG
SHeN+er+HkiZZBlwgRIcEWFUKq+vmb40XLt8gumnwuifU+O/rXsFpJjEV2U+nplaS8+XzCRFDUNi
jtJmCFa76XnvI9EOm8Zy5JKnzNz4WHe4Hzw/gLOW7TStMfFjvExL1A1NMArQHy/ECZD7GUlnk5q2
84RNdMzseuZa3HTeXL43Ku793fCWzegOiFnXJciVu9Soj1gdBcY0NaKVBP/l5X1VGfhplgXkrxwf
g9vCa5li4pzpO9M7vzmbxjc5MtNQlaXsbLS+CIhEAOsu2gykAazE5ItooHvsjXl1loXhVH8BSMFq
OBy1WuYNEIOZ79cQELjN6ocWwllT49qyXZxLcO/clLS0CJpwER/irJOvhfYqT8cJb+QYTCnbCdDO
blZU8o0oTX5n8FG1leROnXZPZ6306qCVBhCQpiDpiGveuJqR68QsZdUSPEEBrYYE+1nID8vsCDZN
n49ePkpkTBbr/sKLbhW5/8RplYKTBQ39/ndgZdqlHcu/KApE4eT4FfffN9FwsB7IznFKMsFvNRGT
gmwJRrOdmDutFsagqZyXqiYJgWaW1+ARuExSyBZTPUygdDwC9RmPtcscj4mJQW9WewJlyGD0+vsC
g2ENjJNQ0QyXCN8vpQ5VDnfrbhXxLYD1yz+BsUijNIp4OSev9J4A4pWhb2PBsDvRcf7LJBNh+q0c
DIdYIf5C3r5oFH9pyz8wHo20rGGYwqdQhaHTtFnvur7qRQ8azGdy5Rx9PlgS+eCevQ94zektAzrB
v7aGWGqnNWqIPtjTkjAJdlknMQmkPZYSDYi0/y6foIrXD1EMNNcY86cVq7EdRvSlwZbsmKjg8CHX
BWAhwWBfgwrtMaJz95ST7NGXBsJ7/9FiPCqPh0gpZ3Q1GMyoQlq6LwA7BH4CQSiA2iJYpodsEs8q
wRhtrS3pANF3Bu8Jt1uSUbjrCg0cTQtyB+Rje42Osz62T4AZ611D/T2SHcQSAXf6Wj+3ze2CSIoW
S+uFif7tmUAKp4XXPOuNMnGC5hgq+nOfi6XxwQOfQ6rzQXucTnMgGfFCHQUyWCyQDVmBMTrGJT2k
81Hs6FKtqcS2TyoZcU8yzfFwdcxf/XTdnT08+5WKElN2QLRFcSO05K3ijVAoY7irgCCyJQWaPcr9
nQR3YAvQ9O8AI59KRT9Z6qBR1tOid/dut0zrCnei6F7rFmCT1Ausx5gml0zsPqel/K13M0/Ddsmp
RE7PcEnmb0aWmHB7x7PWw3b4fZ14D2UU4iKn0pxwpQII8nsLDCTMqINoXnkc5D8pfgbZGVEDtfXJ
+j3nDIQGvsKC3KMDjTBbGisAMYGDAHPNUutUGdZtCnzNXVYfIctIvH69hX8QU1bL4V1vXOTZXg0R
yMf9zluEpRSlpmzkCOWg7R/00wWoCafk0YVHDvGLYYogEQcvZGwaVkeiojLVkmc6zLQvrUI1lPXv
m2UsySk5D/qk2QAZrblmvBnMJ+ffWlegwWpjMg+dMMkKoviif1sPXECytH4t1Hlep/rTgYG4c+5Z
SYFxOyGQkKr1o2o1FLVaOTMiLrH7rfbRwma0FwulimcmfjK5mcwrKrJHwLhjNxiWQvxzwM7V0ui7
B85GkTceZgpus7M16CRDZjyoIFRZjgkufKBX7i+zIlK8SkfYJD3IrzZzvQcXc+8ai+HKBv3V0R9S
F0FcGX0K7JI5DlwlawD0Mr0+GcXhpyACOxtGl3ku11H/GcPgnNsN58tUO/7qjfGtijUUa040YxpE
1awmEjeBSH6wncY+hMjhCozaxodOMh6weeY9cHmwaQ8KRBTO11r7VtFjWgKcnmrAOE1JsCTiWKXm
YFY08laV08MgRgkdEpop9OuWUccau8Thwc5w+cnaKSFzN8X6BiDv2Bn4dekA3Ku797KuOkfYDsfG
6K6XAtoJ+sy0D3LJGRT3KZoasTgiZgVD/lVUQ6OZRYIr1oRrUZQ7zl0A6XxyNkqctnoMIjmyrV/1
KI33N53Lxru9ZAPMhePaUheex1esY8kj+tRkzNJ7jzW4UDQI2hqKnlC5+F/sN+Bf53LzzVwUSR0D
TP+Q2K0S6oj6d4cg6Mr06PrBIOye77n2g6vwMufyRhsJzE2pOnRvczhkOqPqegQI/hhABfIHEwPh
I1VtxQ/nKBxm4gJJIUX9tZUB6yfpkJbQv4FurciMnmuN+MheebpCo2Ma0UHwTt3hny625FbOaA5/
E4Hv+7sJpiYhgAXlSWIUNWhay7vppSnK6zbWIAccKGA1Sx+MVwWtR3su1pf96ZX0BkUk6RxGCtzz
eAWIp53hBMcN29RtGcsza8a4izN1xiIcIU06YaQkrCzA5ZM0iEkDSI8pzNfGCoAThj2LEHM/3i0g
nw/Sgxlh6e8VNP6hTWxHy2u0m/J7OacH1xHyAq4JyK0p5+UH5lTlhF8b2NKYIqky0HLBl4ZiaXNM
NXsteAoOUcKdyehIf0BsSHTJRQirMa6zu5Das5jDmYKvEuTbCNaSW5fvDw6cCIOndq4jsaTVXR5d
tamxNFQqK557wJtIVwpHMzONyLCMjAaX/adEpzPFOyfAfM3wtkJYdbR294TxcoFtqmXqmjgP7vlt
7DXDG9lxF5cZ2wlvQqtm0Xj/5YFmaxnCV4T1gq+CeFtd3S0lGWVJTZ2lZFGj2/JkPHSnPT6SHFsl
zQNoe7RIKPRCYDMHedqQqOPy1M4xFQkGcz2c3DPizGTzHbOJ6qQsbvZnuTTUBPzIJ9oMBUTV6OfC
NbVJE001ebs4vBq9z0qr5YuxK830Ya8eH1bsqof2PQo61mJscClkJWvpKr3PlJJgYCO+P/d6IhqY
Ux+7aH6VB7tEbiKss0AJWVJBwMQo1PfwVCt9I134oNfpg5vmtNo9qonjq1g4L9GqHT3Ye6RZTiAv
dIpfIOpJBpQHWe7NjMVmnuhz6n6vOy2kBG1upqoNv4cjB6nvlHPcHobJs+2U6kJNESQRrTw/T9Wl
RZUmzCpRYrcR1P/9IQLMxayk+KEVfVGlfUsV5HGk9ALFWALbiDz3DTLRGIXZEpqzIuHJU14QkHPx
9lr/pDs3bClD+wMyB9JV9jZPsjn5FbSGTBeF1040xbmyM3glkKopIYWPhL7+uMcVJzJZavVzP2Ts
HOk7TOQ5NWbKjT0fX7/Ymuvi8JfxmChNKcP8qWimWnRtO8yMR7a/bNTo0NOBjEzALGyFhGF7Ik5i
VCSq0ZieszYtdPnnoOgHY901rvypkZA25fv32L/5bALsjmC2C7xJqvr6WM6fBgPAo+/yyCoMSDV4
fUIldkp4dfmkAOUKcNV1gm5iMzc5eWSrH3lgIqbJvh1SjhDGnD71TuLg7knq69v/Y86/jItC4+Sk
J1H5TzA54hyh+TmGzRE589+0xvsLlvZUNzgnnCK+hyK6DDgQ2aka7WlWabg/UUe+QMWcrp06j+7v
jcUjlys+k8ukurH6BiPtelH7rGCbFLhAueNKoJzE6f0e93665dfj0EEeXs/RE83VGduHXb/xjbUz
BNLItfor5XTmPBNomy5VRYV3CyOkaqUP9ogtUeXsfhMwURO25Yli6811uiQY7WEHdytd9dZXITDt
akm9pbJt+nGV/gEsMwlb6iO0YMt7Hm2RLRIfhpr497soR2TcrLJmY6HhwluAAxijrFM96ahAaiiM
iD1eu0SJ/eOQtaFK3XotqcZM0l+X8huvNcWol8A960i7ZgWTtA5tBOOExSqzVQ3Tks6B2jqQdA62
QMndwjuXz/1XBPuztF/JUiPdBLdehwFGt03Qq7Ndg49JWxOOv/TLboAfSO/AA+aFvqzcs84rnD4a
pk4PIJeX2bonSjNEa5LNCSAbORuXmurlGTNGEqxIeBfg3kMl35A/7FF4VHMEzWSv8v0a/sX0E8Fh
Mic/rMV/YO3pOftd1bWGPHQX467gyqoC2JB7/6m0Gr20wXTGztAMGiJ6MGBrXyPk2xabT9iQoGwt
lnW3I53X5Zw0aDsQ0jsxb4cIRD4b9y4a5a0cxrtHSh/g9pru2aub3q+G0C+fm1OlFKf4iiYu/y19
of7kI6QjsMVnD+qamnMqbkN+cxuiP7EeRWu6/+XsUMcZeCgpoMtsxk7H3L2dRHB/XzEyyNNESCg+
wwKFqZDItkytB2vEA3b1aKimQ8KFvthGQrA2OMjOQWhJuANgTCuPHdYkx8WWYy2PzQ8yU7JCLT0q
O18kJmxxRd4SCIb0ciXbKXP5EbYj0u7EU0bz0+ucHJBXk8pkOJcWuIckouniyRFmeo5mLbD46OXn
suwg52Y7AzTIZyOQUdzWJbhtccNb6i21ELb8HfA9misR20In/AY/NDQOtuHbqEttv3dQJLvA9TC4
6TwNxKX03hschRErzMnA7H0L7+hhJ4CJ+g2NBKKEau5jA+wOKviOX+DSZjbBQCHxJWVPidu3VZxb
DlRq+HZycQk2hEP5X2LU26sBjgI1WTO7eEPiQYMHXUxGk5Q+BxrL3FUrjWbO4Ntl4t4InCUddWtF
GCRdcqlsdhIl5xZCwtVanDrE3AvMl5EV2X34UbrUMN8nP1lMoqOusVoUazImoGS4kv3b5f3sUGbC
lmGPehN+MmD9u6gqQGOwtFypTXS28BC54LxXyK3TAdjivoqCxHIVZwAPNWAskH0pNgU6Gkpbw64I
tNcbJtwNKkHfpxYmNKshgfDn5arpYWonInUe6kKPLql7ppnYZyrNMqVquRDrE22zkiWQ1abwktyn
fGG8c/bL8iqXOWISLO0Z0Rk69qKp0Ex1cAe10LSOaMqobfxNvm2aGfvbQHPyX1da7GP0vGZNR7u3
UYpTtOvMva3lFzkSQOsCQCNdMh/wGzuB/z3XVlWutNcIY+78dO0zCbfMpN2H5fTwIAzOHifue+sb
rHIdUXIIJSmFyuJctQmukmtCl8UmqtIb8gq6FDLVurUHCGl1Xo8zjBip65iyFgM/vHvXZQ1Q9ofK
s3L1+uO1h3iVoVTNrQeQJ6sEwLEKI8lFtyEYSp57S1Vdf3BXhbStS2QKJeRYJP2ZZSvA6KsnIzGK
wTfyE8QnMgRa7UXQ6KoleX39OLn2fMH4nvLkzP9YWiONS8SrBtnqWO+gVyejK6zMLRCKPrF7ErzC
r8o8JRh6tBW80ckvozfXwu24bUFk/XN4vs+K1aZEflSTvdDWojky0cNw5bMCxEUNkw5dWoIbQAvB
R80Ln8Jh51LCc7PYmfCPWJ0m4S2Z12VJQ7KJFSeOKBxfoIDvJOfrFMdkSMgS2jTaOPqk5gnKI/D1
K1vqZsqcLNg1IJhZEKwWt0qAd964GolJxp9+RJW9I0kwozh5UhKU+WIfiVZ1FsO11a/jDhqJK4Tq
gJfU0w4Jjzji4lq/jD12t7I+SnFCxoQEvPBcvpRlhKOwKeFR4NH/RtHrdkUicgO5SCqWysHQMv6y
o77Dtd0lEzFrbAHX6Qy2GK0vRr9LSae5V74LrxHSEyv0gxfZ8/oyZECkdE8ZoT/+usxkJe0QF+xb
BFljBUY0ndw8cNgsxMUdKGhyNmPMCdgBOxDWZjnN504w+kZKaPLemez6k4Qw3n5buEhMNI4h0xp5
pHiJ/2ihIv7iAhmWZ4sPcMgcQW/xOmtfE3lirE6wtUrnQT1BEu6pk0zBdQsjh4P3R7K7Vx8ihDk5
PZkdGSrL54mWR90YklVLVlvL065CdTsGWOG+GHW9AB/CC1hW1+winumw6W6q2lOy0kAAxs7BLT7c
UQLm/Maw/G1H4nCMvjG1DZI54S23dXTaXUp3mJiqtl6oQhd1x22IWKxdH11Pa1hhhyoW0Yvknn7b
oRN0ozBMyln7REKeaa1ngZkaTYguLkrtu360OUv4iANehx1TmlsTputth/fCCum8T27ntWYkTcNe
slHFkZy3pXOjWmbfqlzHNpWxruULH9N2BLtcXrNgsIgNP0YcQzq5MpqsCyz7kms/yW2M9xui2cC0
SnXIWHHcA9BqUIlvc/wL8Ow+14qH0Lhmjbogxz3AuByWtsfp/L3Ei34Ik8iXtvspbVTY3miRlzx1
i6553/DjAcSH7QYXXqr7OPrIjSd54aCVjV0VGcWYp1k8hc+hckxdsgLWiTv/hZhx7eRkBDMpKlh3
EezcjRyAC77z1ys/9SYvx0B4D2un93+NGB0UaYr3Ze9mshZ3Ji7r34KJj8mURmvKLunWa8gCRUDb
N0BL2yc0Sl8P7wOc2c2l7mZWbNuncYhQPLIAfLdLI41t2UIBpuccb1YQCuAfmI6tRsUs6iS98oaY
mkB2QIT7fVmLTH5iCt8U2jBdevwKeahvyGkXKqD6+aS54gm9YrssOx8gnF8UcNo3+jnxjPvfqjK7
7D7/czh0gzEhJPQFiHbVdAmMEo4yAlj0kjLxeFfqTGIJGbnR3OwoqGQPp4e1YJwa32zIvZUwA16Y
rxJUWNYy4E2+8dq9M3in8C64Q7EP2+jO6Z5RTDm9VT+skjqQEz3Qvwb4RAN3AFwfez7m4XaELLQW
xbkTM/LrFgZe6wM6MDYgaWjpD6zsr5p0Jn0HEJDYDBPoVOKX4qHpiyM5kVO7xgOMOrT7nUS/9/pn
KWq/UkmsxqXmhMinkgiLe3E70sFofDJg/uoVsBSCZ7bRp2X3hm+4a8UwMDoCN96f3xiQNLQClsuW
I6ICZDOGzalvZPuExr2Idk4hBQXy3v3rTHDHvc5pdpvgAeJG0QPE04IZE9HSiUfLViJHMuNdhm6S
2ErJnOBfHJl4QnOtR1E7txt0scZNJoACMLW3OBVPg+b0WY/nElHvz8RZ9VfHcfRpDBtVAPHnaKUK
zhTCqeP3C/fmO73Kcftb21z2uJz2FCgaLXHgDZY4bZK7CgkYUbWAzCbyWEviUtDSGzL+I19OdYC3
tPDGry6CWzmnCDQ/rHH+w7cFUgGIU7HKbE+r7TTMOf1vpc+J/0iJMbFziYPCwOrsTdGbNwEfsYZH
FabkWRaF037RKAYuV1QUnYhni+Y5Q1NzZyDv6wjPdhLwi5nmofkWAQoRf5dqhVmTSemY/MOSMOC4
AMS+xQeqQUfeV1jGyCq9flh8O8wvAMlRlUAfKnGEllmnqQlp4GqjQg5a/hlrfIWoNP+GUpzUqRC/
KlkffB+83FhJAej+34AnfRLFLd0PwVxz/XKjgsMvongI6YUGoGJSCJlGX136eWL41UUAQ6JFz5fM
v+2R6v2KbN/z55PUiSXuRdYWnUGZNyusN+BXJO6n82UKEMhi+AVyfPLYtp8/Bind4Lj2cA4lYh15
+m9yy+lkzYtFEbQ+zmUp131G7bEZ++PDdsucUPt8vntQfk+eXjXwRF5p40Yjst5485UyRccP+4Gq
GQYKWeThRqUKU3xg5ONgdmBO6a2IqqfupbDs1MiT82xjr9EFgaWolFObhjgHTYKf6Gb6dzXGY51S
sXbXRmuFn8CjCpXeNoNuJiKZnr+9kpRTPcmHuS6fGrOBDaNB3jogD1fk9181CoEkpwrSMP0CRw4N
3/XH/hKjmDNJfLZ9HQLjCTtAOzoHz2+7uc1CfulrcJJIbBdKeBDscgAJmjbEGj4gwnfJ4yjvE7cl
cHE4bVr3txc1fN95N/QCdueMYcoVh0/YUD8g6w7JU0S+mmXOlqjgSbqfZ4jHig5+vcYcjHZQSiFS
VZiIwtsQm9GNmvVhz0E3g8WOvfVuMmadiEE6YiawEqa8QtQzaQnCCd+1/8FuqCcykpuBUVX9ixQg
abPjpVi/aA+jUiK6K2evTAsYJYGA5uDBjnXyg3kyeW3YbYNBpGtcL6p+Lzqa3AFig8pIml7m8csj
EypGisOkDNmW99ost9QdFxgm+D7LF1ur1MjdqwKJkOTO+8kiInlq/Gt7w64EggVyHhs0auI2hOQF
hFlJdv8IurjRdlEPY/uUit01VOWrBYGflNguxHfU7JrWt8rgwjWuLkNmOEYGfCt18j+f9f//BxsA
BD7ipWO7a8iE7z3zGtTWCm4JA4O9AKcIvDk6NY5oUesqoujWkRwOHlmJ8WT7Viv8+V0umE1bcGg5
TkNpB5voqRdqznNtahsZmaEcAVMdNMZWhIrgA1hLmI6nKj0TTc9C+boQl8kUWP0KcBjsWdtCtPLW
aYPdNyMB2BvpOVs9CSGvn7cJwCbk6fzmuV+9bAet7bcKFf/jiV5f8jmmc4RTowliIHj88ujsPDED
5Zl/x3MABKd+yVPock59JkNzAOIl8zlXH12vrnDXN83VqeGoGbBCXkl9YrA/Hq6022Ses967YO1N
GVS3ss5KONJum9YfVPgm+5pyGHpK5tyqN+qFJlZept6UWZlUJlnInLGKUrmIjYlYGVQAljlBu0ZY
6XaE7TueIDyGRiUgGJ72lDqkK00rCWLoxvwMPdinSLdnKvOWY5QG9IBwJINw+tTNwCRuBbF1Qawc
TRTT7Jr8nwn/gfPc8ciVQANOjDVZrTYoKiNovy5Rqui6D3L9VawUbJx9u97eCSVIzIlTS1qnHxOY
vNDfgTXIDX2tX7wwMdxD108IsKpOfuFLx3H7GYqxBlRon2uOGbB0l3RIVWAnqKPKfhj+DhBg9cBN
OElrDIztLrLgHVPtXBK/ix/t9xj/E4qcQE3OdOZc8mXpBAut76LX086KjkI/Ag2N+QdQU1MLKg9n
qUhlw356vp2cJbJ6iS4kQQc4N0ppEHnmXPFJt6sHy27vU6f3Mpl21XfGFtRhjG78svKfretgBpn7
7UmbCRL9M0eM+PTopUDfRNZ+BNhMt005V2Pi/HwnVw8FSuGcdXrX4d/tXnnYhr1/cUr1qNbc8PTy
2CRjXwsPipZZVyOsBL6uA/lUbnBH6GhaX6JNK2phIZvhLryTcdR7VOGW1p/LWpkN4/Uh1xdPzIoa
/3JQlrShVU8VFcAYe5uC3YXsXIxfb8o7VUvkuzvlgiOaQChPgdca7g3eaW57944WUJYwKXySd7TA
C61yvF2hg1150GxGHz9f9FuQiokrD4f+Vc/c4xk9+DUonPmEiaUA7GNpRgXZAfbTTnFVkjytl5qu
/lD0Nz6I47jZ5MUpZ/ACsJqo0jBdrNYSVuzbZGfOyMF/FnqIGyOVA1WLa1EIUD7+ENw29cLGkZ+g
i2Xu5zyD9cAqNhk3Pam4KeV31v5CTmxFHARL0JKyw9fNlK6XtwKoiFBY6SqwVOgH0nnRNVTYE7wf
WXibok+ahXn/wJUuGny81FiCcUJiONRKKXvY6kiuvD9bzYXIUnDNR/IzraTKYwoOuwDpXc6mq8Go
fhir3/vmDt5xCuDlH+xa8ITusuzkoYYTn5GHuyAU0KoTgiWZUlJH1oGP4m0yk9ivfC9bQ3NYj9Xh
U3jnrXoR+dDOaqSnVpQsBOOIJ6iHNZSzg6jjEedhCzQOVJuhb5hUzXxLhz1K8uVsQ9fdXwz2J6Nx
13e5PvwfEz6/Hda9Ebbcf4CGTdh/oC6VUY4WwCIqdMVJAWx8xArLz2hef/rqNfdGIPAEIGdHWMMf
eoLB2Cx8PsyrIIvFqAe32FaG+xKBMS1IPr1IDFsraIpMbBJNnmD2Y1x2TtqyVvl+gef66mvbyt8J
hvMyhGeYtXHDec1GEXGRj04ymym4+4RKJ+wuL20aMWSvgONSCJd8iCVO19TO2pWGAgi1ZO/qSyU0
bIlMsGhSSVkIumsG++GeRw32MySWVcRvilYjsA3SbMc0S6YGYIHROreQbBzBa5yGr0fdMa36Xr3t
SH62j/tBy4jxKUbsryfmeuFPYYz41Grq8ZHeDk3M1AEJV0U/45eZx6DEz8LwCZSUlMy3XZzGmFuG
e0vHY2wNhATfcJJIFB7PQpXTFiXvHMbMpo3Fc4UY1nWmgJy9AMF6uX8U3G73bPMcgiPhusMuFgQT
Dc1rbBh7kgenJZMc+gM/xM1LvMub5I9KkEAD33GqmJ/I5fWlGMGCGK4iEaxFk2WvRMQYGHfu5PXp
ulOcYb8O3uFAJse/D1pdrs1g/mNNqWWgyrO8CYsZR2mJAvcU7nlTfpafr86QTE54vq3sa3M4ynap
z9oBv3+b/c7PIAupPIiwjYlfW2fS3BtUnQNoxO8jX8OMKjSHowZxRy8JMT29uIJeSBAO8irlnmas
HT9sdNcitXU7uDMqMOwueL2j3mYPMY2tJg7Z6p+CkV+jD9REqkWVl7W+Z0uOqvJUO4NIWMazcc9F
/rR2OaOT0M04/otX1rWtrm7DRrkv+WQWrJUEwDVWhxyz4syJj88EG9KjUxh9HGZ1iODJpx3Xy2Mf
mLYOdThuBgBR0VmmJ+77CUyQkaMUuSEU1TxoF1FnVXffWYVCj/Rczv67egMT/oZNHpiDP512GoRF
KTe7JvdRYLi8s+MG8drx8PKHb2YXBHItdu15Z7HuLdyRJs27/UmI+SBqXRuXX6dRUqJXQP/QHkXC
wKe3A9Zj8l7Y3cPoPg7AdkwCH4DABUhcxTu8QYY1m2OvFP/i0jsQvO6AWWEg92ccm0BCseunHBlB
sdYkgxGz0mKV7cPfriDucsQAOijH5Br0LeqEtr+ODhSLKorQFKtBZFnLcm+02wVHhi9gXTtkKuUo
Pbi2oHMt2MBPQgW3qxSiBOOaYjaqZ3qsrUPuj15CnAlOwT5VahvTFPI8I4958z4xIaAyo9ZBovkl
zbIQr/1/j2fhYjgsZZZStvash/gf8HyKomjvta7o3PILxGZpd/y/NCwD6gKchR0r1KS9Pm0YHaWG
zK/fv8CIrqVRUtgIpmTKL9T7i8gMcJEVh4USdYHuqnxZSNH4k/3q0Z1lXkVmeQgxFCVxqhIPoZYY
dyydTsMhC18QJPcdp4Mm2Z3Guhj9ig6hv85d2fjNwbIGm8QxY+1s7RKyImx6+P5yEj/h60NQ4QiW
WgOrvxHlUvtVgJqMuZH2NRD2tzimKRUUWMjWa9Bkm0cPe/AywISAa21gjQhKnzvYncB5tnl6Isn2
zutMRS09hrw2FJPnWQMwdQrhJz6oYv/I17ReeYm+LJeg9WXFv2iH1WmN0Mg7eb82ls6OnzY4MVkT
R9cTdu6xW25CNPeildKQWnjb195dCkQ4J2zTy65O0k3hcN6PoWeIcmk7DnmWeqtY39NZvgxpD0LR
p0mOPy7zlNYc9baWCKh72bW3ff0pENATcjpSnDhtQJj0yOYZV2DJdjJC6Fe7V8JSow7t5Io1t1hm
zFjak+oZxihams+Xono42QomwBfqoU1p3CJmHEoIzrc9kHqt07l4VbEFHGLV6ejLmd1gmytCj5s/
ZRUuLESRzd515a6/axqRSOCQ5h6DetMm3/PO51rhuqaBjw2CQqH2L4nv5UbUQ0/TCFdNQzF8xE20
Kyo4e8lgBwIv0RH2c8gwGQmOOrbjQWr86j7Cy8u0ksE5Lwg+GxRUcaYno4HqHIfhwoM4YR7QCuTq
R2WjgTkroiZ5d5x7L6b+5ty26ZWKfojH8NG9y40b1I6L8FIZrgkFrLuujekSPWiD06FKae6vTFHc
3lcTPvvVYBceh5Ik0UI7cQjM2fYCnGQGWRWhh75a+gofq5JlbYTeMjSLYUN3TxIF3p2v+0LzYNif
MbFYlo3myusGsYPob/Bxa1Df8WwsDeiyAakalKu555pkFbrXhiPdrJWQ28won/eKrwHTjYLLiwjo
t3piTxA4ESeIl+3O6TE4iGxqTqgH+ytGs6ZRcq5wPDa/3VazjFVGIW7R96c1PYdpp33KFw86PXFT
a2qF9rIY9CZwRfCNLlYk2/NvcBynWqv/1nRmtIQcEW3+dnPGtZjio6kU0cLGHx+GhE9O2PD4LBE3
8pM/64D1xuThI+zymouTUsz9nbqtthwTiYUO5NG8SWe1zXaeE6ik7M62KI4oipYnNiLf9k8epdCU
rwLgNsGc8RE5qyTkYy8F03bxOALkxW1B4TCLpQcErTEEIdnFPUJGNwSsZVO6l86bpTtY/Y8u7Ni7
HFCQPU0msdaxanl/GdPNRHk7SZ2LSh0yK0fkhdvBwzp0mBngrIJoBJaRCjccIKVQIXWDP86f9dsm
OkImjHPys5YdG6kh/qspvAzu6k5xpibf63Vvq6bmHL96KzRxS6DAzG/Me5BSvfzBcvt518GBXsW5
nxYAcgGy6Ezxam/9oIavzGF562FsinxgHjbQjfEB1xiR2mG+uZfmS67sXyXMNPb/TmYouYG8O31P
8jH30dsFrLqzSM8EGR4/uCwd+58scltzLUvlngn0QWe2nbZ18qFbJbN/2Q7vp3qVJNcwZrBoonVZ
j7FKcmnEgVAixSax4gb6pSNZYHnplr07NNgAetDwa7SsC1BtuF8sLZLTACMHpx9M1fAbzDiV+1aB
KkQXMA6UmfFaYipwcbDSnoPfDfrbvWF6Qp589bPT82zGJMp3dkx1ORF5XWWrbmvTJONwMu2ZskP+
pohQrnaBr1IltomoEYVN+W7J3FeujlOt7JWuQiA4LL75AxIhuoN6ing1ka0L2eHnkH/5YArVEYUG
eq3FV4GFQ/1/XaddobP6/TVXvW1t9PRiq0Dw0CVdYsU4REtkIkZSYm9cX7lNO7Zc75Z0QcyrSax5
HjrPwEiSCGPkNNx42IFEaQSUSq1Xf7FOLjLZXX8j3EbJZG24pP4pBien7QEPbFe2tdk2H8thwgmI
ljSO+DZHOFY0AWzgmp+Q2kbpHur0pgUB7rjERr9P07d/zOZ+TnvR6cBchfgilcDddLEJVxa9zjV+
ea5Aj65ju/0LQpMgi1e1iCC7Fz8fPtyQwvkba0H86X3TzrWWvE+RwQPc+8/sSKXuRKC+JbkZRXic
B5EVituEFNvrl4j1aPTxyPxY59kDiZ4oz+s+vK7fhRp6LhSLqjYDE/EmSruyuZQaa6+nofvmt2SL
tOQ6g+6Dd1WONp7bg5rZaelgWueGoVS0Tnu0Igp5jnRhP99YONZEdpNrPrUPEIgHDo9m6p5ideu5
LF+Mv4V6pcKLQo585ZYzEQS8JTSYOJODXg7StitLVP+iB2bxB23e1onJ3pD+1X8XeiohQRF9JsFq
lQqfWrGCqq9x5M8qZmbCZ+SCFoeMadPaxGdMnjmwaqwVAURYYjSKjKsxt9L+LRdsYCrlOEDrJYa8
sFngdVU3o3gaKiCkQ9prFyJa+Ga3hfgy5RQMf5/UFm5xSNUlUtVIeYPfbIGNdf4vsPRDXoY81Frv
hCIdpmBYAr0WHqGj7smLwnEyqSqmYwb6VciRJNJn1dGj8DIi40qh0vvU4HJmpngJDvfOteDAkc5N
Qgr3irZ1X39D2XN7eWkiW9OZz3gXHCUgBj2D7xLSjyWVZ5d5T5TKB1SCqkHLF0lz1e08iXLgTxCH
I+zHSIPEEwBPWdyfPBcxGG1IX1qG9ItMmC0Vwgt4g4XF+YRQe5BMiFD8i8Xt175vsZ7cBSnT/f95
4nZZKNOEc+zPO3W4zk9qhKDS1hLIvoTItGVR022KFgIBuJO7Ek0+zLDkXr455cqtbsTNywMno53Q
g9U6PzL/ycgqI5r2Oj4LqPsXXHyKdeDjJpd5bpvhgt+auThTnPnuZO2V3XlOWtU7dRCZAm1racFe
FhR5lh0E6MZCi46WQCiKscVYRYOMelSJUgBe/xGJdVZdeAnFTEhvvuXK3V/fPWoFlKp27VzsXfxC
EID5YrqYgU+YyZMYm4X7fc7qKs6nbRAN8OAWcUDpZddgBTNsfkXyyUiB9/lqmYONZ3EAERXy+Jd0
3uQsoVMUaw0yPzIuuo1Cekve6qPQYVbGGEUqOnRbVFQx5O7MloGB7PdifTpmEM7e/d6XzTSedc22
leXVgxcZML5ei5REziXBy4++g+NJjjWRc7oFo+q0BDTAymGRRVwdsdWbXPlkTD81E9Dg385L0Lta
WAxt/WNGjOYVxYwSn//wbkit1QeqwamKtQtsrefzSfJT4vjLvMVph7iDcN5hXPBpTY3gLW6nkWfp
bhVwcz+NF4K3uoS0uLpom4dvx6hGEdP3U7yjqEcf0Lq/zs9O9huksji8hI39SrJa3SuHkP2OpoD+
fLe05awijFmO0Dk1nC2MxsH2jVuvHeVEM11Qrj4PV/jS+P8ckdS7XOc1OecGYPCQO3ipz1DU+1rr
Q+4vRpRWAxxMSAh2joJ/FNqLyZ8P+fcavA3Fpo5wx1l65JaFfA04vpKbqA6pLkrpw9dDVOWz26WX
PMb65J6MTQ/umNjLb5s4Gag7CzWPeLvM4wBgTKjNf67dIpiFrFVbjQOK7cv78OVZe0/SBwcUMiXV
WZrvbkSFPnjOLw/6Lef5diPOmdLH5rfORe1yLW90CEYyW45oIov0572R/0unM0J9nHHlW+ZlZd92
qFdtWWXFiy783F4oPOQhEBBBn5iFy38yZkZh2TaotXJyQ78lnd7JJbcx4bm9gijqv11SaW+L4yoI
ApoMowyzHN6MT5WnIINdGEljekgwsQLtnFVqvELVC166jLwGw4NlrwvwOo6AvfhFd6KyJli/2h4p
m0En2KeJ+rWUMWvTt+1yfa4Ux8suTVB6kCBStyllvuSQfthIAHvo4/1xsNgga23lHXlSPPqFrB+e
ifF3RX9WV9NvyE53XL33mbeiy70kEEi9lcRlcltLvTvhw2T+SpfRAHs9wj1MSc+vFEEbiyZ5y0QM
TkbAHmcUC6HFlOyIzbARLBBEvUtOS6BrTb7tz/v1DwSXL3FApBKbh/DnpxbGj8S27EGG4Vd065C5
e50G+Zcj5m59/bOSHu/mnL0I6be5t7/qc9CT3Jh9UhA9jxmCAtWF0Kvl4kygheOE737ybDHHmkF5
inr/nBSMJ+8IQ2RqUyYYrhj48xRkoWTyeTc9V/07+CkYt/ACQww54A7ObtbYzTzWmDqaaIS+VIOf
ziSRAfujDXGRK/q3L881bgd2Gr8ql0wZJnD7FSLs3IEoFSNOBxfP26sKLEPMULIQnGMctHCfTgZE
YdIOYUBt7s6hyBIL11EtlSHK8PkeoHDxAw+unrDmQ0bGR3dHrzvlsXd6y+JwG0vnzGd9ZXJU73X7
IfqgYx1v0gfMXw8vjGU0Kp9dJconUFFkBByPhb2BKGhGlP5AF8G1UIWchquH9IaxJ6Iu1WYSmDnt
pjP98ySc3nTEmHvQeL14hi8hkdfDU6yu1BmZnP2Oc8tID+pPoYsLJ/bv5EDeeZO5Wmna2w0vaPXa
nwp7/8LgfzRuQq9cdReuOdm/fuEbER0etdsI2XbKzzDE4PpZfyga2ltAMNB+iKGKfZmVOVjDvqNE
lcqUPRUm/5annKYOoa0NIcBZSHzwFKdxgff6sJuUnaNewIKpfJ1h9bNIlP6tE9YRhJRl0OZZsol4
wi7udHlBL/W9Z+LkoDDHwoxIWkNmeCoa6TZm/KX4DW/eIqFYUJJ0IJ0YScmTcz16RWY2AO5iDQNY
LFJmB8XCd45AUMs2UpZ9wjXa36y0gvIxbyDrU/DKwYGEpo+HsZVxfU8UYjXBjGeuO4MSuOK3HVCa
5T8eZdr7jKcXw/BoW2k+wRK9BuyAp/9VZLot0jEHRumsMEqZlxXCM4LWwk7VXAWQaTrD5cL1M29F
5N+uR/8p+zlYcZ5w+diQAkzdL79ZFTODbf8tJQFVY7B8gkVLaHyHy67nuk4lFCvgsDmxhe7HO16Z
9WXdbBcQUc2V5aiT6QPmv8zXBKG6UXSNDnMiN3T9s0XMR4yMJl9FXE48n2HyBRNq56hG6kb34WNo
Cg6MSEvqD8I5ADFYyajS72xDg2kwk+4WGyKzaz04bdABvf6xyw0tx3HbYTL5BXvbwp4qaw1Q4Iiw
OkfEXh2YliSANvT3bgUEATJpFGUuo+5Owr8kv9KMMFR2GGWfLTsT0DYJXhaA3x8w3uHp6z5huFMQ
6WEawaKWascjrGgrIB9tuoWCR/oMkYCjOV40HyPgMV8OyZJa12znrPR5g0EzD268+TbLn3I3rfgC
6BnlUnvOAJo7Yn5yvPSlKsGQYVNhCljlaTGbxCxkRqNLbJB3AHNKZcry8Jkk38WKrmKfaSXp32KT
E+vMhk0V5j2k58MLVLQxRtpadKyatG8eD58klX36+D5IRW+rhmXMHHLdhsBmvQAN6PfMJesYWeO8
qIWZkfXXd698rBekuifYx9yBShAtPBWhLUqvhtZuw9w/wkvcJ48pE0GXjsGEXvoT+8Wz4cMikQ9v
p7Gtls7yG6igg3dqzkBNgzctE/sW0+2DpiSEl3BhJWZuCi7i4n3w6Ch312nxuLTqpsGVQKZAseqg
63UIiy8bZE7boH6MZ8e2vX8ZdzpHss9DsNH50NbLtI2+rqsGjKk/HYdOu/kqE0HR7lhkiE7HmZV/
5GktJpw6RBudcP7EqO81PdY4thlqfb5PxZJU4edXYkWKET62mhfqRFUK10N5nCFXoxy7FNP+ov1M
h3Q5vqUYywsnfx20sYSy/K0q8KT9uRXEsZ3QTo4mT6/JIEM3+upT5uF4eu0wQQehDN91nnXBUtZG
oDdcRC6cG5EBrpoaaWsLCFFYlB2VR3xXXeacFvIofAmEG/CVlGHuxI9FmaHKOXU1zEo08b4gINJ5
je2pfTRjSQhS82EeKoM+JlYGJjxum5Or7GHB0Ga6P9E01URbNu7gJ3H5lvt5iIUMWY3NTSAoSUSf
Kc76gRtV2LISRTFT2lgpAtGecSE77h2CwSiEh1mJ3nUVMDDQj7x5gJ0fxXldoh5+MW+5l4x0N68o
0EdhqMOmktyYoO36nHEvack3mAGil+lyA8sFOrd0oHkcSkqeGJiAqBsBu4PciXgPbMy7OiVERhDY
FjQll39eSRKKN2Ufv15nWZCfrdDIu97xeY876beEhisFm1nqFf4SfQMe5Dgi9iFip11XUwXpHzJ8
MYuPIEOYXuHHruj2wUG5UIHZ9QhY8ovYiTgGO1QPc1fBo5N+8VvQ+LxmsCSsVcRh+XavEwgA1LlY
pORcB1GVBowkOF7nMAU6jA9B9MtxtaxRoEMvkH3R7AxSW2PRZrZlsLpEQtI6LDiuBvaz2jdJpeo5
f8RZtvmCS3VATpKS5gGONzZi0wN6TIebARvG3jGdgcQImneCOEsfm3Lq17BA5+s2WnI44avaVVlp
oavzGwdkXGj1sucpt0k965/oPK8WyV8Qsk8nCnH2gY/kyrAJLBWWxzwoIF4zvYYPVJmOADAGCfJb
CVCLUNNhpXse9XnpHYhiDFnWtLsvZtLqOTctJE4hx0S8Uoe2On7G40iE+oargsZncjToL9zdEERk
rqYS2jA8xlmrqQAwCdw+nHeI8ITl3DtkCoj3EIBPgHfYn8hZZDm4VZF+9B9QWzq7VOJ+0SYeFtFG
tzhFuctK5ofhJvUeD81JqB4MtJC/1NAgptsh6+qW8NWCk+wenyN8KPLtKG5KJIwAK4rW6SevUHvT
r/qb0LAB1kuIJdlSRLBSlo6/f29LXg3QKDn+qSEQpyShj+lRi4FFV2MB+zTCWtVDt+pDLu4qPlBI
DWuaQ37c+BKn/eeDdUa7bfjexSe0WdatSTygjoPMQ6GaOcARaIMRhKn4b1zZ6uK+0xRDdprgpIlM
9KH6kXhWTZAUlOododnKLSGYCBQn7Cxw0FUbhm/IGqlX8V+b463BRJHfpwNIakAnUBdic41HWbQv
MXNh66vy/up2vyM7jIZC89s/I1OswDhc+OJBNcqoGZ5rvpcZLLcXrRGCI2rcHwGjCfroBThEvCOR
vsdn7TyCZc/dqpi3R6+XIEihDIa6ms91jAPC/Mu9TFAh9wamhvk33LeZ/TyhiOEzVhHLCnYICN2i
ZabzyporWsqThQCVblGidiaf4pQMqQoZdZoY1F0r3TXnwdQrFmEfWhSqM6ktgoXwWkyD4jqNgZcQ
oxE20L1GRMxmi6X/AxZUbAIVtaQhicQTzgNacyd4SyDNUDJOK/fQZOMUlxC7Xr1wrbxkuaDSKbxk
h+3+KRBcubL8JHcHLzziuImj8bogyYeE4ip8/mk0MoRTi4uYfYzXebd1TbvIybbU6KpNUCGzvpy3
VryvkrS2YjAK67YJKmRQIVvsdDpWnmI3IZwgVtUtHm1q+bsMABTiCg/D0JE1HnTlLfuUqp4vqVxI
S6hDmVfxAswl2SBOq19RelmhAasZUJ3VXxheVXdvQ/2IiSZx+lJaPoCql7EAoFE+sRjskD2YhCYe
56jPMbLorvYz2+91y04WERvITDJ+cJN7JM5QXdRkO5UoUWeiNJwPLwyGxET/01p1tcRAay1ovM9o
bO8CIGMihn26zmFsmKl35e7HioWrd457eXAaXyQxJj6anM1O0Z7eHGe6Xp2qz4VuRdPwG05yFuv1
W2zIGa7Gb4rICeUDdyuvSGaLM3te81ZeQO3b7S/sC/SDFDLfZJg4nT9XXpPvtgh2FHG2PaUufabn
5Ia47SbvJn40LY+vXH79QngwmYw59lVEfObBFTI0vpGs45knAXf4dndMBLtD61j6aE2pJHGlaj8a
PwQBK4dWUhgSEdrzow4pjy1kD/kRNUNw6fNKVaNj9j7LuzsAVXh8Y5CfCxg/+5LFWpXC8UrzXUXG
5trA8gI7AA0Dg1/3uNzxso2CUljUw5Ku2S9jhSHLPTIbWxOmKQfmEPRaQ5+ulSV/2RsAbP4H8UEU
aNOMM8NOottTq/bKMCrh1tqLadJzrcr1WtNbgCwri6fskQZQufjKZxmKHAC9U/jZP4aMcoz6t7BN
v0695kngLJ7pNyin9YGhr1gVpQgsiCzh2EvNhv3bXOd0nVIDZLSRc0m8I8EswhS3xk+mU44R/nCK
SoprHhEAWsi7bVGXVS/Va1bDB8UrMKr1fb1OoTvLcUTb8t9DFhSubqwd8BM22+u/c9mFP7iv3rEr
pe9ks0yIXOOGRcJ5/f5i1RXZLUqdMA1Udes1DvfsruK1E1BSTYx9Tm7Y+WhPo1Kbg5+Xo92K6IaU
2v1+PrNug5ZzlyTACtHfHfAR2pagvJJ5GkYnCGl4hzfx6C1w/p7y9WTyofA31KSlT8wIHoCXiF9z
/TFvCGeWS+A5h9auVUG1fbqJVjHSUBLE5KgurTpnhLt3Z1fQsyLKzDZvmFZ+B8QfIMFMiaMQ7mpz
xz4ZM5r4kGSVWCp9YypTY32MPLEPCHTrgCibgqyeqeeSZFKrRWiWZBC4C3vKD9z9DW+BQLdsHq5u
63S3oc+hvVXJArt2kjFwtHneJqEhsdXLLTDmX4QiQ7TCLYfPf40YV9EZAF/1eRVMO9fatXJM2+9O
h2DV+7F5yeFxZdA8Ms7jsUSuy69/nRJTVvCCYjEg2MUFHCcem8Kq0ywpdAk1bJ12OZQ5koR2NZJ7
yiUgasq5IhhNvcjiwq80PUgE5pnoAGrbbNFg+Rqi29JAenuk3exMTI8rCWmXitnTsF/7Zwf3oxan
DNuZ2blkCQ3q6CVZMC6a90oDePQvlBbmvIXQJQO1qI+bgOvaXOiVEEmbtR6naZei5XcrJRpFNOpJ
msUKzu0J5AoJ5SLy9qox0E6HsJ9uxHQlJKFVzp//xf1QQVrb3FYR3iLD+tJV0JR/cldhd/w4K4p3
8zPYlbGQaXF/5/LBry3/UniYSH57uZJuSQWaN2OdT61//jptwcDnmSavHJ//HxJXYtdD45J/1Qqw
IXs04vyYPjJtlsUFU/b/Tka+dxTMMkUM0zWuqWe7JiGfCEow8aJZW3q1KWk8s4lprSEQ716y5ULX
io+wOEGIK9pR7KbWlNs3Nt5hAQKzTcOVgDMWRuAEUmGdYviaJCCA8QA8eHG8ma0tafPu7SoFHV1X
vAv3k833dUwd3undCq3/e1TdQJXDVE/rZ+BP55NDWL/Q4iMiEPCwfn/N59be1+J93TcCN+d4B9iQ
dLAZ04gCyXZdQVjLeFKbOjezY0pPmEul8JNrfeCETVd0iFPdfCllskiQhXOmUmIaE9YLX+fGWaT8
bpOuJ+OoQ6z+NHUnXtL/+zAe/axKs8VqGaLVEuvwPrCeQsSC8hH9TxIWSkzkBvNhfqcUn4sx4mHQ
yxSbaIutocrpvpSZdJDqwpT7xRHSNESGRR5x2fRPCBCgQLS0ilMnEcg3Q0DpOFSfmGNHLwOV56Oj
d+AzCnyFAQAJdTsL9vy6hhcD9FzA9MleqOsXqowjmJjCdve74S7KycFWbyXxzZiHAavi8J0dPTn0
oLTyFekaPr9JzWlRyh3Ad7s+94YXaYygLcCLdDY1l+0xAw3iAjch0jKkXbmAT8ZEG6Sy4SPV/GVN
g3FnAKqywb171psolGrJ6Irty8rBtXp/RM+e7Nz3NvcOAU6ul+hHDNVGqPBR3JKJw2um6j/gU0Dp
3nLFbzdKqvQ7GXi9cmQ8ZGm6rh7ontF57SoYnl4dFr8VooCXyhpIuwtbd7ZsAv2UmNJ3V/6UEYwH
bXFBbNeFcmhnC/XK/myYT9cqHL2aWobNq4l4bo8+/GO5eAyqPkdLy2F9bNqiYBeJyn+XBfRL1i5/
qVggrEuyCYYXZZnAyz+T8U47JLuzQi3vkL+SOwb2BNu9Rl/ADRbD5PsgneHYo52DWcVj9pumW8YT
v4Ujno8F5RdveDAA+NhATUQlRSXFL1/QK85Uy3VYsdOskvym1nRpTcxThFY/kBRvEdOubIVisSHd
wf0t66B2sVVNJu47Or1pLMrRhDW4d8yJ7ND+rsLu7FXD0Cu5QlVWF39DN41Kn6N7UwpPGc7A0jT6
nCE9Pwx+Pd1tv7IXVD9Yv0Z98dDCL1ffvu2rapF0ZSmmsYTeE9+H5nCnsP0DAlHith1gKTfUVIyR
YCtzqEltx1K0RhECYzxAg2TpsYddNZIDhg+9sHK6LUk6Xxacqw1n/7ZSpIfDc3vldMoDkr/hvbky
j4E59eBuspb/PHI/wOTA6qcC8Prnwm7eLJdX1S1rfAvZnVS8mml4MzUl0f4fvyBWvPrakmAWMniB
KLbe/L8AYffRnPQpNVnOQl3/aQESzghfnpF92g3wPnH2tcBTsizerxsz/7lHhlmm9Ohyq+BlTJx0
AxsuFfASTl/d6PzPquDc9n/+GIk/qScbql5n3aBRTsYXTlTwmrHtpo+wFu9zjWQBxjax+Is7RT+Y
VLnMLwH0efYl74s/wFICLcWGR0XiTfmYCbl83g+m18ANr5a7kE6sIi2RuQyferTSmLE/rhiiVZbA
f0THZWQMRN+N/7wLUy3yA0OdtrdrkrVGjPomWJ1L2KFYzlQZiNtiDodp6ygB2kCsJG9j+KBy80lW
WzrtYgtBv5zbUhqnXkV6nQTuVdQTj7qKtBc+bYhhuagjt+gvOOjw5+wM3LS+vc3Qw66fjpen9Z26
rtHcpoNmV8XhX2XVeGllHhk2zNtvjN+7Bpoe9idYiq0YWrVe01LDuMYU+rdpeogcnZbI6rtEd4aL
uLmJBDMx652Jy/4eZY8M+7S7KBYXsItH4VKqjXpD426rT0GkU5LXH3OxXajv/EN0eUCYJI0rtDO+
Wok6QkQ581MV2NWxrqxyj0zbGKUEoK8t9hdK1Jty7ZLD4XOXceErzAJ8Jsgo7ZDsUqjo7fbEq1tp
JIhA8ks2AvQy8BtvEZrYRa+flZmxN/EdV0dWEnb+GnJz+iDlHkSvGHnXD1w3AID3/yBSh3/+gMx2
ArBrMOasTeGIuOaZx/QUrPMVomXog6mdeQZ/61YARPDB9pPpvkJbivMWnqAu3Z/VcUNnkQ/serC/
/NW1jZEEhWJjxrTZ2yLl+Gzz/DcbBVTeB1FHAY7ehYg0nZ+VoBihtmJgfdzcC1FESImbD8iVzqVy
7xPKPqsxzUcwM4Z8wzXECcvNMZA4Oj0b0JacWON1AxxSj6ZN1+Pb58A6LA0BFDC1cWkWPUXbhcy9
d3F3qxIgauAPt/wejdDitNg+5MOTYQWHsl4kOjDteHqIePuSPipm9UkFxS/Q1STHSVtYdvKjxA33
OBZpx7x4w+p1L1mVTwOPurDgdbmsONcs/UJNovWjChHk82sYLDMjJiMp6C1tNS+3WQ8OTK/27XGL
sr3cxV+fiuvjzs4HtidknxWWj2IlLyl4TZ2Su39AV4iuM82lP92dvt0xBucBhXDRvRbkr9GeMemC
u+LvXjy/0VGqKmbIx20aXD1GX4dhCzgVrsu92tgghlGOuJyWkuXkocLwKLjCAWX12PDL+FuIpnOG
1SE9LIas1Y8AQMVP0CPwJBbQgiXNDXXX/G+SyoaCYzvwbco4r9lxin5wN4f75y4IngFHfXG66U8x
KUEqSAKi6SjnMuqhBb3DrAblvgEwN4BnGj7p7U2S39DQxQEYS32ouon/IV5JR0c0O0pEPT22PWy6
jfEIEM+VTd1wWmiW89iSbde4habkBNhnOr0nPHt19x3/fTR1CcMyd/GgHw+ExQpgfU+PgDl3Zq6o
AANGH6QVyCEdxr3zLUns1QNaLIGmZjQMF3gG8sBdMuqQP6iHZ59zpB5Bs0EwNrRkwtWJpjkjaBel
vcFbfJnSbnF/wduxYTMmjGAjt5ncZvUGXU3FxXZdMsJAAP158eO2J/jQTUL8e+yaw5GnTLIJDI4M
h6inqzNJrW0f74YusyevDjYv9gDfpG3tGu5911eBe+8ymdkJwIKakCbDAwcmS1ePSBjOtboKqk9z
bAKZg2r8HLMQhWW1KfHlzivBteZubTvTMPTWw3iW55fws/jt2jl+ZCIidmPQ+SuK/wTiqthreQEe
Md67V78a3nLN1h/qq42ucUULoxttO9DTaT9FLvxvcA/SL0fnfWX2UBKOG2sIPLoDfRAW/eRzdACF
X55gcOMmIYwo1Icji/83hQuPHLfydgNcTijrhLjfeqPUwC2+fOBWGV5KkZOk15hhdbMIQqPHdwoe
7zhvgtrxwkq1+vDEDfcYvNS6Xq70L1fxo4Xzu+lIT4L1yU/D0VdbQTWW9aC4el/CDAFknXccSHnU
3kdsisjsw4fezA/2wLS2SfIvvCUj35qYahjm4V9MXaqqsBBCKkZKB0WUPKYSn6f8dhBwyGwdNrV9
49tQIOm7B7dopDBLgua7Txo+HEHoMiSqcdCh7hXUKxIdYCdzYhAX/HAR9htANNwb2LdjyCAZpecm
SWNfkOH1xBiWTNG4ChHLvoqIuUh+ja+opIhl9d2VLAH1UkaPUXi8o9Z2B3k6WEoL3+yBtYTN4lfm
rvkuuSNFgSF1F6R6R7LxzeUMbwYB/lHjO4scSOpcMTXx3ul/6aMHhDJ4506VboXFMUGWbRTSRan7
Kjk8pYis5B24y+2oqfchtVkJh6myach6v7Eq13UyXKx3mBmhXLBt4qKcpN38JTwE4uliiaB2986G
LqH7U/PdmGdLkb7QKXX1TyjJavRe6YLVjyUZIERYapxhb+AAFAQBcKjGO9E8By+O7m6kecik9Vdt
uapqnhsKVoVkP6Itt5lnpy5XY28R4k699nkep0fwau70B5wog14c+d5ITR0C7Iv2RgA+3TXO2Ris
hUneuw3qQzVG53RORH+7JqDaIdVCinevV5kuFwSKIHykFkYSrnl8v4xklZY1n3ghUACZ3Ubd2xPc
QTELs0B/H9nt9P2axcN1+fYxEufG3bA5iQns298gwaKe3xF+oKkYkZjxuYEefX2oF0K1leuszxkK
wpw93JL7gSKbEhcT7lQZbSbKBMorhfhnxR3CMK/KrtoRvLY9cn5PWzJHaFtWq4bPr866XNXFG6H/
MeNrxUDPhXuUc4Mf/qM4Qnij1FF1+PnOYEu6DLWn0ERJOav1TaBj2mzkGK41PpvkU+0N7iFMxjir
rL+YxLgkF9FunjFQ/vMJO3nnDHp6FsiTc4L31dX5T00bNJp0U85g4crYIpnHeaW1LeVQR2Jqzjhe
omGZhiIP84S5tKoRwRaWLYo/Ktkgx6Kk4QSCDaOfrmH/4DMyi+wNoHw+bSDiI8uVIQcscajD6M1F
gZj/lYGfNx1YMCshoKIEJWwUO8n5tIsjCZ8bprZOJb9nPMVepqBrkUdCXH5b9AOxazovzBdk/y0v
czzXHYoCXcKiJrcJZPQhT70WaP03a+gL5M1OBKQ/Ws60OzL5LI7WbHQK6KfgJcGvgNZPoQISdkoa
xyFEJRjYrWUZMK4mUqQ02GjgIExUyfEvISkcf4e7h6Ns0Jl3eRU6xct0QyO0rcSm58Cdeu41303P
7PnQORBRaaOh/eTvYnxLYADBu1f8Do3NY+RCc0NA47uPu7RHkOwKtp7Ly6Qhb7d5DFyV0/Zaunkm
mCKuoV9IS8SM24gwy4Cnlfr7u4b8SIAS85VoMI6Raiti4JUfH3UZJKPyeR8l9FxINO4IhQZurM+B
POQIK1YINCHAKeljc3OYPy787YfboC1i6bA+wmba4m/GfcgbsNuYS3bC+llK3yYtYll+kSZSc4hg
iceyewgwHoRzePSi/8CMbp+FGCFRaPQhfUki6Z8n9d77Hr8mcdHooGjmy5CTFYDBxO5EdB//sdub
qxnZaamlc1bnt72zhZmvR0HspnayfL3r/0mbApK467Lc0iWdUQykjMgYG2u2SLxXuFhKpeDyhJSm
sNH2OYhg/dHbySIekl9tf7DUwDD9544qbss1Lqo1T6Uxkl8Tcnt84jubAfQ3dzq/oR9BgCTY4FsH
YKAcqwbgTuNE6F3semjPAcbBy2NHNr66wF+3J/aJEytichQNYKucVKXcTzk1I7XfRNeoKHxzr+bt
bWO7GSaP6UbdtKyi8oFC/10viXdYkkzCr2kC4IjTtzKgcEEpbdP+3pzV3bNnU6jU0Tta2wBLb9uM
LIFeOyDeurOF3UIuCDNFXfUxMCAwUiMGxiSzMHZG7MY0DY4rc7Ue2o/bABnCjKWg8gUEEX4VUyzh
toWeyewVmiGkC3MY/3+B4Rdk/UAFFQiHW8aUVXqdDCN3hqIi7og2sMR3eRN3V23ryISdaFBWVA/c
hQQtrgTpkmwL6mh+qhkS4Kf4f6eoFgJuQvAX9uSWCwmZtn3bRVSn4RxSXRAgSaClXiirTYsa5ZDW
OAYzomvTDJDIncH0MC00PCBdEKT8/ytQaTKyPQNvnHiuKWUHoH5DdTHInD6EXpA0LrnY2EaoC8Ll
gKFeG6ZIcncEJlrsDU3cxMFYXVv0DrinNBHjibSSKklB5qgMo8Z7W0pdaBgh2TyemYD/4+wSt5vO
GJ6eGHI8CEh3UZe6/NM9gqxQ6IuXNn6BFVZXFxx4/OWUmF1mZvM1SIRsRXdvvTvNOPAuat7c9HJH
wDY/Y0OsKSfP/UOp5XLiKW16aRLF2KgHorpz4QRwsNNm+IrEZuqbEpWhNJIGBtYynPE/5ekrQJe8
MUgwpA9NjBMS4MOfQ/7aXg86CIApq6HaWVB/+H+RS3TgtiSjOFB4cUhPhnmQ5+1+BNWHmuxC3ina
beYdTRfnaLjfOkuTitlwux3x6JxQawAtjSdVGFF90amWv/zfkDsrFcDjjs7e5mGlKhSp7fjIja2k
a3C6M8D97TYP/nyMm/oOPiOLgvmiCspMfh0e9E7urisTMQNpzEu+zWRGlCNejxBciIOyhLZA5ukY
KPTA6jDaee13QSqOboiuw+E7bqi57KtN1YyTCxyZ8V5XsaYCMbB/sMF/+y7iGve7BkslB6nAoHrk
4R6L/BZZzyxRRwEQz72h1OmgLtBzd+A+d6oBsiUUpZE011j+DiRQb1U8CEQdewjrGVPRRzl1+Agr
+gFyjw57GrpAVDLAc14CzHFutzuHCHAQIBSMIHRICoNWRYrmZmpDZkJkoT02RuzsgrcsmPRPQw4F
9dP+Ss4jvplRPO/lTJk1AV3KNfLxjf6eTRiNnZltkg4on4Kc2xcD9ZLbawgiDDHtpqYVFBmXyHH1
wBemhB+PwkJ9CKQfta7mcFd3U7AAWca7+CMKZe/MDlyiCfIEhK2VPhhu+aHpMnPfcjRNQESPsr33
oXitLQsudg7icBWn0jUU6Z7+r52fNqgmLk0ifIc2qSvf+rksMwZ5TBHGnLW97pBnuf09psIUDDAq
OAOTfqCoC4M/70yF7WXbekHQ6XHlo6laAvka+e9y2DFE5rCaSmTs/3hk9xraymfqx5Vau5j/yq7V
rvoqvM+ZmcQct7JB2po9PFwWAVWI0Sx0du6FALbHbvJyKot9ERhxTYQfHKvIxhMuInQHIoMkBOfL
EmCj4vhc6x+8a1rn0KgptO1KRoNjak2kJpTxVxg5wl54mqnrfOExb9AcVjgBSHjrzvAMIJaokrQy
pmAnfOj6o7xQnW10yN8CEA+OqVF61CbAduSWH6UhIU2DSKfOe080KSpdFNipl62fh9llXbg8/Z9D
LBbnx1GK8zxMmIqpDrCfJe7Umhz+JRbXQk0nEnaMdU+Y0R1T9StSXOMZrSRQ39EHUu1H5S0BmeOY
pF6oJNiUc6BtSfuBSQVxrCOlzoEtE2R6mNPLzg6r+ij20OBX+JU8N7bDmgXbpODmW1zbTcZPe4FB
xULgNuNS1CZyUmZGlYH7d/9F+QNpbygMLKlAgj963U9aqJQ+as27JHxxtFK+UFDrfSC3ypCUUAE5
BDBQFo1/Qn132XMDRxq/6XVvkwvgxKCqiWMTW+x5lJj1j5XUqMBTiYDsTUBLWTvRFMojtqFDe6Oc
v/W4m6QbkTF/1kWvImHQpICikeVZsznkIIrWVvTEZ0iKLdQq/M372yYHYqXouf8rSVzaQJyujeva
zVrIxHfNU2pB9ZJ9HL47jobUuiaH3ix9/wG7MrguwXRjEIJYqMOWpHlChaJQP30HuMzo/RL/636u
OqbtyQ5+VNnL0bnSgfBTZrGXpFMPdIBg73H/uPA2JP40YiTvLqwYfIudo0K6H8TEKXCuRZ9PZZ+K
/tzpZDeuLNpQNWVjPi443F98pfrqZyucGZz/HXclX5ETx1YSKeRh3pWNM9sEbd+W9JVftP1jdhec
jW8LHZaO8R1otnrORA9eXbv8wZSPfDjBxL5/Z/iLXAJqSZFfU974CpL5MzZOK4xhcdglU5pPkdL5
pSsb5dIHFn36z7/rt9AtjDC0BLq8VC05hXbjG0gpNngInpEaKT1057XOAyM4RPQlDE/WW1cX7wfy
901dZHOcMz++spO4C5l4h2FBwFw5q/NsdO7Z8+UO/2yQuxszNeAdO7Eio8IjburCz6nGWNZ2MLbZ
0oCaBUx4KtPTslEKwSqnWPuv74aY2YCiibNLqmLZY4K18ewJeQHuPKAOfhDaLcMT2eN8Dwd1InAZ
xq8Fyj6kDNepHses5PbFtWwr5K/d5zvJmWeHHwjZscB4TjXjuR7V8Nu0PgJRIKUw4RJfDn0nZu4D
cLdX6goAF10d6V/8z0IZCZwfuH/x+oBF6Xuocbk6NOdwBaZnFMmVpRnoAFvyncnZ5189F9P46F4h
29Kg3oLXc7ROgO3/QmO8THVg7qKI79VVJSJUUNG0NY8whowTZGfDv5Q6fhVNeMQrxMtl/3QJWo/c
55fe0KFfTR0o0TNhtm/Ymzg+mQJzcJEbLXMSO24hRmO6TpkfqKI1AbLZgLj2JZY+wnlF1qLvXSN1
SNoc9au6S9QwXIWM9oDBdFJXiK8iftDNoF66p4YT6YxokXLQO5sSwKNmMBocgdeW2zM6JwqWZX+x
yh+20ACW8mraYYLhapSmmY/Q0AziG4X6oRDfCaTlO+JUT4WYueti6aISftnLe9oWbb82LXrNovJq
ZemLxLkSDSPD8FJHM+DL+zi52RhNrY9xbRRwJbPOKhLdQkVVQJVSf32nHu1GOriVh99cvnd4Zkym
E9G5K/X18z7bD3WbqJMXS2CGYIY4yVLtuX5eBOMClgkGwP7J9qLAwncqxdK88X+vSgoGgFeloUKc
RIZcECzatPoAUM/KXEgYjOZbaTenAnF1ws+IioKURqq3mAeVVgfviErASn1h87XbgfeLok7IdZcs
ZXbqJERcH+aLDe1Q8wQqKp57xqrCk20mV4yAeZ5R4eaFQ3ZnCWvUMbi15mAQ2sLg78h2w5Zmur2M
aLX/fy5AMEE0v7bBsPDO5tREiqedCMcrhwjxUHCP0v+0SnntVOox9Y83O5Qsu+vazq+3rM8vbJP9
FHddXpPdvw1nHvHNiJ59EDjHC8BEm5Z0BmtA4geuUpmDjq8NNnOu0xjDZqX6aU35XfSr3Tk+UozW
XVZKpprqSMONrX0VzsZdggdKXgtIgj42+YQSCcEA8luoLLLZWOh7Ctmr704WOZsnPpeDkIDi7zJ+
MpXDuIJUeG+iGDiiS6reWA9bB46psHh+E9kPNhD2ptWHN3GfOgvMpbIsWD+s70Vhpx1w3zMtmHa5
htakr6igwWI0zBQHM068lQG0L6pZMXVdRU3z+fk/gI09frIB8u9sULOCCv0qY95r+1FKNCIG5mHH
M/qdGbojiKdWljsG8iN1YYmsFD/QcNNmCWklxR6wAXcGUTpRDQCn2tqpfK6E8VRTRJ9H6aF+3W6B
MuMhGxknZ5316aYyYSTn8pyOw2UpUTERcXfQBKS4MFj/JK6HaQXs4He+OX7nOn7EEjj/YEZso+5x
s6fclxr+ReHSJswJ5HBURivL7sjxsrAbTXLkCqFL2/kV+ZWEXl/lI2XHsOo4H4Pjv3v7Plm1qa2I
x1ZRry2HDuLCcLO2Lp/ehWmscPYlLeiUsqtzPP/3H2XrL/QYdxD7y9EIK9jwQrZusSlgEzw8R43l
hJ4P96LbjLCM7QEsuNVld/RGPyfxn1yOErdqYS5Kov5md1Cabmpsm3/F5kpeqjokN0zvvpVJ51z7
hlLeZkKYTE060cLMYXDH3CGjAp15ozCAYU20UZs84Cz2QpZa9C62EPy4/kZj4XWfbxo9+rWlNmrE
wUXZbV7RYZVdKf6mAdYYInEPNwx86XIrTsgB39gt1V+8O8KXbLSf+TwD79qsCa09UK/QpYRQPKkC
PBQz42aDbNxPJ/9m438vLtjMolN8ei0bHIxSQvTB/gegunV+OrlNhD1NbQVUnsnPiMiL9FJHsiKz
3s3u03iriQd4zBpmkk0DJ6G8FQlYm5MStR+MlLfgD7kObb2/qMVMyjj9vGrUXMgs5WBRiuLorqhT
OcBkDJR28JvCvas9uaTJTIzNGPe6mz2s+JAhGMZEL+JPR8lVWw9SxtDhRa0gIMeC5nuzwrEI3WQ1
XF3z1dIbFB35DzhWDcHqiatooXkn5RCLuN+Pa/ieVudb2Zn4SMlBhYxTXQa68fcl7blVkfMK+Ggq
xI3H0bIGgsrrwQdhLDvKWx+KDgmBtvoMSLhKJyc8Ht4mE9oiX8ZB7xsiVXtQIQtSgUDo5ynS6dH9
ZxLd0E3U2cJ7DcXqec9IMJvinYp5RQwqjIAdVNKBV8V0iKM6cevoKjsDADztty7W1VtfTUTrmkUo
YFcEgTiav7cncx8GQqDTQV0m9GjCKCiE4doOGqLM265Yep4l28Id8ctL0N8wPQbA5hlMz1Oj79cU
LH+9MkiHSWYH2+ZfK+p10Lf4g/Rh7yusQDxAiqO3x3Ow4H8CQZHjnQcZJGbLE+8DTuZgIg46Pd8r
3utb/j/4MRNNVVeDq5gr3FN05CSspfm+rBf69R8uKIJXjL9G4xpFkmLFa3lGyq1dtN09FCYfqN7f
Hx968XA41mZ01iDcOSOEldPCufMPKx1iRwDS2RjIvum40bYt2/oUPcfo3x4HOCPh8YglQ0xali9/
kaLT7940SfH76ndQTHwWSjQSYUM/usFQrZIFBrPebUKQz47XJsLNWUTagmlDdFE4f4OG8yHpu/tK
S53sEi+Rrb3UJqAyHJIvMPBszQdJ3k8hQNSm1JgYxJHXm+DZX43Enh5+Ganq5hD+ARrK29MOybDm
n6UGuhOiOCnf/BU6llF3JwYNqZoJobGE6cvgJok0JBd3xIm7ihSzp3GhA/F2RAFyruGV1xkkJUNx
atyTj2CyiLGVJ2P91bSdHT6RP/oAWtx9NlVUpyzhi3BJsZiQqS5LzLcRuyHEDn5tAsTQ5R0b3/u0
cvv6r4+1xYYLLZAhzo1cUb+6MNB0rBayhDdOUtRcymjdJxBgMJXvElayzuuFN3GLIl7vJrj1uRaN
pgVozcWO9J/Ico5QtFxPRm5BWayUiz4FQNWX3RGEviimJZ3zfTfbUd1G289kTfFnMqq8Yb0yMRfg
LFqw27tPXr4vX0xq14yD/YsxATdbHe0EP+bKpvhLB61dkyfIRNJFevBxpUhxb2BO2kr+r4JjWiwj
MtXVN7STxb8xDRW4haWiRWic1mp7jeG+kUDlyT3BftxKYPoqDd/Sl3pnHbqhzQFefmfo5yeFpWwW
h6e+BcbxKHw0m0TneuTKX2Uq0FKrw07FSx6ijJos+5H5bfUUIHwEbdIksu2xHr8dM9L14ENXnQwO
vevaei5uKuLx9ErY7nRBoQD9Pf1cpI4Fmwd2lWU/AFmfENg5BGUuoEFdO1QYmElm/0nXZoc1R1jU
JqtW5cHsIudTH8/Ck4KogRKqX/3my141xqpdfZDh6IMHXua3MA0iUvNxZWjQKTEUQNAWsEWU+q3f
chiHzL2oJ537LusX/YQ/A9dYq+3x/kxEN3Fzwzt2q1HB9AnJ8P4vvbgF5SqhVm6Uzr7sZ1vLaR5c
pAW0xP68S4NGQgInjEWPx/JKWqvQ5rGZ8e/KgwNb/o0bupTrc6TmA6lgeyUy6mfPypd/2Mz+gTkR
rsgyx0eM0jZI+2tRSNZUUeOpKcJ84JBn0TnDqmCKGj3SlfbiIyxwLev+xq79bGgj6XNDaId+RXNB
e8hXvktdai2sIhwFUAGs5WI+mHtaGU2IBHXaLL1bN3HCODyUsO4/15VE5YtjrTVnVfOJWhfCfmER
nlObXTdAMN8d5Kt1hbQV8vlo62k8NZ1YdZckk0Go6dOn2jmE5vjchnecioYSwCfgVy7i1LF7y5xh
YEy8XK9aM0uJLeDQN55E6rwrexDGVhwHGHlXfgDrK6682ZBJN/lzI4q3QbkEQENZf4T9TgyPLc+P
GrECxmFKpVQKXuPkCTGm7w/xt1Yc+7Tt56VDRmsEjcWHMo48J6Tra9kpiKwxKxMnqhnDyX7JUOMB
DYUAjI32Bx13HFC7RTIjbSv/x819ObRm81tPq55hF4iXhR7SRQB6LBaAJsL7Bqrk+WdBATkAiRCQ
2UH4v78J2abGOFya5Pu7j6+bNTLRcixvj5ePxtPhzX4zWVcCH4adre7hftRd8tzzgqPzFLhibfFF
jP/Dy/ASJL6ZRoAWIjrSS9L+1wR67n1LNgxamR+WK5nndMgjcC/eJrQwHwV5iBR3CHbfizVDSI0u
f57ACNwebPFnY3p+m+JvakcGunoK0aC+x+2DQDg2MYEKDQ+DJpoGEwoAMmfCD7PKv7qyDw7hy6ER
Su3TvLrDwpdynv/H1XKUo7Mi9f8qWYMWfWY8oz2csfVV9RbivIxo/AjaiSLGyTZw9zPl082u7vpR
Yt3ZDLuxnqlDrM17zCJm/693ufGl7+K4B5073lilcFtqS+dNsASTGv/EmbskW5n9nuddy1r8dKS4
HkSMSj6YeOKrbUNcYIZN5cghxfMsqW0DEtgBQDuHqzp7N1xTn2OQ8IGrdntFg9ovmhOvjECsxGME
ptSztujatEgMu1lup5XkG4DIr1IEA/Vod1I3rl+mUH3TozyNtsT45Sse2VND3aA7ywz/J4WffIOU
cl+0a9cpHio7q7p89sy76hVsI8sBgqqoT2ZhSwzvYE5e0/fQmLQxE2oUfhQzWMCPF/JrDUx9t4cw
VrDLGILa0XVU9tQ+R4aHkxngoQejElrNznvr7a8TKhcJemuSL1dF8/goRDYWz46wYJY/6J+kHIL1
ZVJCQD//imC9NOYM9Q0OB6CWxnq8+XnJpuEIhm4BJPFg8PBi7ZJq2SD3Rwyy2ExvvTBx3ijtFWA1
g2sjAsuBATWJKgOVW8RI4cYDkXN65/MLFlW+d7F9I17DWbljFWK+cHHGLIsH32RmWPLdfNffW/uz
m0yntVBZ+PQazsYouRNTSeOHWkjgbPbQa8mmxZOeuUrv114CK+iWAWKkdn/ajx40tF1Ngeko2U8y
tWrkl2qJMRiVCF0ILPWqvD1tDz778W/9sXNLR0gUbY/wqWFHpuZEwpKio7vA6MjgTuc+uWJnvcSn
FNxMOEs9uw3he8IhdCTWiqLGWXZv4ivz+Qi6a51MuATaOoAJpFBh2MDu5XXwrPSc8Ais6ogTfXbr
fw4MPFl4po+B+FYeGm7DPwhvd/mmR9qcKK5Fwn+6n/wjwTcALMAD13fD0AQbjpoACEWRhzDQaHt4
7U85y1W8aIUuGDqCd0xOimhJ837U3BKILdfXcUI3aoyJjVpJK80EFXht7rN0zThwJMwhPgoRb6ar
YzESUuggfJ9kVs14dEd1DQEsg4yDjnp6guJzQtotfjuRh/f2EG1gy79RmzwxPa4xMHaJU/WvucaZ
wJ3Ni1B3K23hHfjQFooHheo5caLjkJ8v2wrz9ROS902tuEjgWJ9cgxZbt51vqLPSf7y0E3NfdTyo
vBQ/EwdAGJ/c01Yf0HznMumHz/8Ikijl8TRM4GFTnDCOn9nplAXK7OtjUxnkebeNM4pOVtDhtD66
lVlJkKm6KrRgEXa1Pu8SuHFNNTETGgF1hc9StVJSNthOf+X3ciFpIC5Uj830dBKVquQhcI37G7h5
XBccG4alM+0wpVoPbJ/yqiNRGvsUkFWGHd6VreziNPZmHqpXxLCDGWgz5T3BwztiYKODIMufEOSm
RoZHSlWnuWCkh7O3p0OgHIfAcsfy/oNt/XpLNbQ6Q1VeRINhRol9iY+4EebwKZO0TkLUeygfd6c7
cIFmKoUCJBCuFj91etjSVlqqKWQvPDktVo0NiuJq2vHvngF4sItsAGWicoHhdpo/6unO8iDoNdvp
hYKBve0C70CrQ81GsEiAW0p0t35iGBxqn0trl/OdMPbVlmz37f5RUT47xeHQtzAgz+JSdXb0z07W
jXKKN7MAGBWyA8dXVCPAUi5pU+MpN96P/J7n9WgrgjAdu46MJkDsF1n8fFiiXpWBmvUpOSYCagPH
Ip81QBq1czI0oW/TlFUx3OlJgvrxgStTmcuPjTBtl6XHdLzIiD2kkONa0L4795NqnfqEYmyfp8ky
zfnN04kI0BVIvam80VFFxUgWlrk2SKkqZXW25Lv/l23UIomEMykUHl/hvQ7dl4hEUCg3SPFzNiM+
U47BjXErg5Xj1B1bike+pHOAFnc9azE9UWT+csMUAhvR7YRWgtTO9Lcd66jTJBp/T5I/mp8s4E11
nU846vU7uYLVmEuElHcpIZAAgJiUcfNSye/LjDTM1JDiMoUN8N6CZuQyQgqBFzHWbHPjkNn24YYi
5FdXS5ZCEEbVUCRL6ppIOHVQRitwAjNtfXyZCczulDjGTxNr5Bp+Z3GDPObYKkvymMdt8nkilecw
at1a2hSo24xgWlMnrjTou54LHAoWE7/7b4JsEWPndStUqy+GzneiQSh3FGHjZa8p/cNilhtF8d2d
19h59vk/hvMugQkB3EI7qShTitEYCF1atAdn2NE487DZyHR4HZUW817xW/ir37Nqb8EjD684UBYq
kE3ppEYxELLqWqvAKkWWNnlTX0CWqeGtGEMS+ioIOMb72MQj6B9oFWBoJvCs4evn5ouXhuFclsUz
I1MNhch0xxRn8zBk+eqN9Jmt3eCi/obtj9KWpyKSlX9YKpUuEcYGiRViYaRtm+fcXqqdtUJqiw2F
jfrNoLjz7XbP9H3kj3bYnvhkXaaycW3jBITFItGKRItnxjZyjwNQvoGEZmSqzIBuTLM8lgOhORZS
0Cy6YtqhPijIRnep+AXZJCVIbGifGN+Wwi+eHIyB0I6m/JwjmJ/+jN8keVQg6M/+xAvqwGfJVJqk
1SO7siq9E2e5kU0TiiJP1C9bZpjE0QUJ/KUzKLS284Xdj2BsUFO14pM8gx+vgfYnIs194yPDahBq
okj3DoOBK+vG2HVcvQR9NHb+15PVUTlz7iWiUT9bZJCzxdpIy3dYuztDU40/pMm6WGjYnt4t5b7u
1F98dpS/vtm7NicC9zetlPsryGRWOwofeaJ3qJnCc9N37ycNK+/iF9BPplk8a3CmtDHLsCMSiVgG
fd4h2U2foUr7uQriaUVu49Ak0h+C29MUO3b7FW17JerYq32Yn11aXsTMbl4PSNa0T/l2Vihu4XC1
eBF/ku+7FfDizUAdIyquNH3kYhyzL2vpLIBFAVIZX97Yqod+hsS//CVJmiTzCQbhvLZlhpopR26D
zVILtsX6TYH7faelgS0Sbdw9G/FAUqHEak1iS32UVYo3nGh2i2JUxpmvGXcPBIm1iEKY7ZI/nwuG
BPS5qTfBp0sCsXJawE159ObnS8LAPhq8SkqaWRK1Z0ukZlu74O/CRTyxcWGfuIwBQKzeqK8d7rCb
o23rPx/KknCLHkjdTsJnbVl8yl2FONV/pMkaGUx7/bsqiU+w7bLgCYCdQvp7S5+ZjvzWyF8AxmWG
PQvayDg0Wi/+iBjaoWFP9CbUXC+Q2h74DLcA6V89VWnRbO/i7LCC8JUwvSo0Uha+AQnk/u8ijS3c
YUEvfCsKR0faMpBN2tGvACt15cQ5tnvV+ENfSXRmqzbpNChD71OGOcKKppIYW3sRrTErCsAWkhd8
7rNYsZqpQxNf6YaszaM6w4Q3bf0IQQngy2m/hofBK3jPdxieXpzhdlvUDp2vRFMUwiNPSXeLNLA+
qT67pVxo3GRbQONa5nnVCPlQ3R8F03Nc1HBTdHMiASbcA/959WWMCFwLfO2u4MSBoDMKTHqu3jqg
vZG4wPfZ8x3LMkWueX6+t6NsxGC3fdvJyHoXoXQNWHiCg0U9ePeaerLOcxkv8ole68Vk8t/LqH8T
tFHoRUeGwJcV8kHr592d1yGEcOYZEuXL4QXnlIqckMQyhbSEEW8MTpovFZulzIdQPoEQ46iReXsr
mrhnXsFOvMeF14+pXF81DbrzFAlq2y+l3Kj3Taa/3VdBl7khPdvzlVw7deMFCyPTcCgaj3BI5vVQ
o7rn13uiBY3159lbe+gCCzywSIMcWKc4pPDtLsxoWS4rzjqKDWW7DCCoIBcu57B8qXEg8Eu/9jdN
qb9HK3Lbt8tKVPBH6cCjQwTLrLI/v5+aTN3GP+nrOj+YnmYcVJjLJi9I+A8805iMCMwye7dmsIoz
qcCZjvVbqCxCXe2sy8+gZSb5VOm8BEYHL7yjOIoBjtYwiFA8JD8FOEcGW+LCUCafaeujpgE+qlXq
g/2Oic+uKkJs3mxRkWzgDzceiymHdm3TSPShSgbYixu6mnfDXLs64h4ePBDHFfaF1hiib1PBAwgD
bq77+ZL2FKyx9qASKXCHSVja668cLZU7KfSLaBNwTYJRGncMTH1u3h5OUdNC2Qc13guD4j16md4Z
jAY1PwAyK1ickPvi3acR2Jud97Ghte51bixBAyIL5jcUZtw3c2fTaRufHvOTwdK1bVL3O5JQzDWd
puat5skZNKtwEw7Vse7jYdu9rdAsFWAFJsD112xBOhH8lPqagCTXlT0n52nc2fEzlXDW3D79Mwkh
L5+upmLcDnOPpSh4kNK3uLFD+tkCxQXRj2p7aHoW2pJuoiddkUXAS6ZVJA2M9wKLfIGHTWNYvPvt
JH9iB9lmktBlsg2bxSc51hNnU1zU/E5+Op86B2Xx8oQaaJuvJUggVgY57K01T1rFykuK/ornr+T1
egFhVOrWBxyKLNQY8u/ITBTD3+k7PPHCMwpvUrQMehAmn1RLBMJEp+sWhGFJURmzXwSWxfOVcxUk
BTylMkCPdo5lTkbkuwZ57ihY53K5R8XCPFedbZvo8giWUEbpRgSyLA97T8H/aMCSfpPkJbMQC224
90Zf/bfhHDu/IMo5q7j7OXlSp5mM29yrlOAdNztejSC+dw9hHz/bWTzRTTEVA7R8OeBmffm7DSRI
5XDFbKnpaOZ/Vaqi7q8+717WJk9EYCvfp5sU3tOVOJG0qMJfXemZPpI5mNGKXnBUkxsrc9TM9zkb
tdAGGp9RKLFa95OVXlx/Cd8WeULZhjoF2Sq+wIAD/li0XKBG0o55Qy7k0ZKKZfuorDlMXyFwTx6I
AWkYrabnKCCm1ESQYXDcDinVwkneW5+39idEBDQSMLBPtoJ4KJKA+pjb7dYVce+qF8/5vHzxpx2d
6Ou4lURgaLRKggOdDqquktKyRIeGbMrVeSbw4pLhZQlqhnKMAIefbzbJHQsSCZ58w7AhJV2EG8Pi
7nYQoUxyRZTnBnCfN3YFDFEgo8OZDuAHw4fDcTFYtvZY+DhE4b+26QScecyOq0vT0glGYeRzRk+e
akDDjI2Aq/jjQxiPH6Qtwq887uiG9ynyhG/IbUc8dvS7BrZsDC9NHAucFvGTUUo5GcjyfltI5IsP
mMcPfZ+D2UExor5eFPLEeALPMzTVWfDBVQOi9Rxv2iLgHZRRz0ixlluuEMEBc+MMS08m6UDwQzNK
ZJagk3CsXiNmXhdqiQgJbb3vF/iBP0fcQm+f46BlnsCXNCWss6mgUJeuD1QX6nXc13WHhszK9mS3
Bm+gsNf6XtHFO0/vQOcv1usPUE/DgeethSYwvGapwS7exThVQ8d2xsXUvRoyFoTdfZp30muK5IXD
7u2H6gRq3gztL+sEYCc4PZLlv+wLt8Cq6ofiQ2U+QWrlJPauOQ6EFbe4eF0cvboHEajhDG6kVpH1
uBoLli1YoGk2sj/932PU1+23rdzNLBAQmRqeBrYFC8+FiuHWIFadYQKEXOVCzITSzGPiKB9jXOPr
EnOlpZKghJXhIuOrczAq+NpYSnmKLzySOZ/z1lhuRXZWYJUXJuc7hLe8Ivjdaz2mpHkonXzsImoU
6B0aN9mG+0QOuxzqICTEDIPrnzXbuNgTSBXfzyrWRMljh3RscNRkTm9xUQB/VuDsYn4K/aXC3pjr
RGDR2ZU+A8QPCAjGUB1iAmIKdoMPrUcC8e3/06yp1cUopz5H6uvt+3W2MkUBUUUzagCA94+wfBtr
FSqIfe3uQPQa8qerMIa5tI7eeD3WJWwaG46Q8tmWLoXGzAMWLizF6H2IN9nJd65fChNqpmv5qGWL
eNOhn6+pycKpecvBIccsoPoRq95l8YxueM+goIJGpNr3eL9m86GzwKR/3GXhsChTLRgcpwygLjiT
WEm+vB2KfKZhcTbXbbUcXbFrKCPmmMB7UTfD3FlYZoSiIXRJft4q51LuvnqIAwzDeB3XPvE/fxSk
q031HoMpSr0Hy4r+zYaDOz4VCte/C3Bqd8FuLLlQmTnvf97DN3MJZfD4R6TxD1U+gol8RnCJ2F3o
qz7jq+gDOzyxHjISVTte2szAWwnXiz91JmaRG97jbg1DdOBfXt5/LngfWpnY5UnEwQrxkikK2DEK
F7OJZUdIIfVBTBJGNQFVgg1WqbRLu9ncO4+EZWYtdkQBovPeskomazZ6wZOvWGMrY02dkXidkfRI
vS92Bz3wIbuSa/kLckTa66lJ9KMtQCiThRs5XXEfrT5aMMWcUyzHwfVmzSbs/JChBrcFgK91Dty9
IVQVbLH774um1BGU3wLG4zofsiPCCj4LFIvFnGejU0BYVO3/wuWYN92LUz2rdH2SffMwVfz/QNSe
CUOkZbcRO6i1r0wBPlSdgoowC9wCbrx8/7k9B4oY7qk/FFZQbx8UFvSU4bHdrG+x9Kgzuf1gkcdC
3qoMfFi1TzG4u/7IktR6/PHNfrgp8pXT/YfP7/8ydh6avooGVoFIdN480+bdidfTPu7bmZyvGRpm
DUEefc0F/3LaHOHuLSTWitWZiUe5JHtvW5od2I2+drSgx/IiATLYkV+YVbNh5f1yX8uSC69qItiA
19JZmsjX4TvIlIAnuWeLzDv57ffGvzSTlIUX+43N/Mo6RpTVcwc3Na7C59lkLASWpMoKQ0172f5z
/GbwwCRTyKPn7nO6z8JkRAtOfo/6eWx5YsUN/aQXfSwck/bAGjYYzRO11pWjgHT9HxHMBnWXm3cr
qJfY5P6uWIpYEeNWpZejEaBTOrekfU5p4XHblvd4pstFhOaVHP0Gt/IeDiYGlamqgnU/MelCbs3c
Z1DBxQG10ITFeQEMR6s2JV17j9n9HEpjuCPmAbJGtKdyI9jk7GGZEFpUsEm5L3e0QDLYnaXfIkaL
MyxGjf9ZLqxrjtWc99pduNZ++Gcd43dztOPPan+eRiUQzfUhnWzoG0XQKyrBKb3kaE2wT7X/ZaF7
PFr8GCeQPWFC84wCg3jeCC+W5UfCjBfSVnRnmQDdK0JvhHBLGLMlSYcohu+9I1R3V9iqMco2xgGH
NwXupaBWiORs5+8CaMr+UypSRWnr3pGsbaXWHFm2gTmB7TXVyyJX0SiPOhSYGID/bO9tAKTUpC6Q
M085+7laKDxlxO8TlXRaNJlaNwBU5YQzzoMRLVkOu1GM6T3PHIM0OFEHGc2BDGFmeoosag3miBO1
KCpGLq5n6FFWXABd61U4gCbUubOK9iocRbuBtFt1KjQ0hIBDkguQhaI5jnEaCpj8DVm88F9Z1d0z
qbfnKCGo34Eo3j2e8XL/U/Mt7660Ddy7MlG9byaBGS+6y4vhPhv4Kw11qjdxBwqxftFCjeRu5qpi
/kcZRH1gnYe3lkmC0yRttMFY59ho5Z9gmKFoKZ71eTIZcZ72jlKw4Z76r8SZrrZG3cQBNRO2eXog
CJJjUmu0ica7jamVZ8jnF0dVjHK3Kq2yRMIZDOQhwx7AbvwnNRy6ICNEhbO2qIlbVAMS+AadYQFo
bibbQxr7Es2VRY4g20ZftSAAhrcT131c6edIJGcf8HuYOPEawUsKLgWodsqI04B1O3kU9oF+XRZ5
5sDQY/6iTHzYE06uoMbxhp3gjrybIu9poUDXa002VWVANvUQH/vRzQaXUgjQPACd7imh6jylakhz
N5tHZDs+5PU+kLEFWA/sObNXBzyiqfsli49eeKlf3aJVpBgyA59zPWDUmJQzt/FFYP76JN0VWRLY
25xTFGP6N27tFydVYnJmdHGfCF/lxgR0nfrAjde3XT0pPK3EOdWFZFZSQPP43B5lpe7AEymSWL9a
8dPZuzkHpuDDx3jZB7i9DP1whzNgT9mw/j3vo7531BnP2TZ9ZgG5QWIArC0kIKZf21ZSU/EDPPBZ
ydNw8gtr26u5Fw1lkt+Bt5cbl3F8MlVRE9d6GaXZEH8CvPJOmUsh+eN327s5p0bexNQZ5Rbdp/Tm
spS/q5sSR1kqGj3ps3XRs8d2EIq5mH8jbjWk4X0+Gxb3w4uAsGmf8+DO/HOZmOUha3KyM0VKKDRf
doKHl+6MPsqOuxU0sBjsUPtTXRZEseHHitM28FPJuBWi6EaoweUd0Zn/+v7Uv+GywmBC2r3Cqb5T
9vkL+S34f0zBDl+rMOGydyTSeM+yhEd/6UY2nEF41YHV6TjUWq4F7YynToXTgzIH9x+Q+zeOYINX
K6zevvo6ppxt6l+ZMpIAlqTCayXk+6ZBh2IQJdRdQ4+blItyeoY+uY/jt/pIxyPJsajVRUWQBC2v
CHrXxyDfYA4cy4ershgkEvYmAVmQU5LAIFYcRlpWlOB4EAhUHsMZW9qVnDjA1W8QKQCkmI9euWmq
/+KajgAPnmt2g8VAK+avpSlbr0D9d7hYpH0HqO6fk/HmqU5f2CBxuQbTTIOOq5ntDXMI6ubs8yAF
9MjxjB80o7U36D6tzZE9YuUqRrnnCUi20x3FW5LkgrUbIRF17ubAY2+bmzuVM6gLEgJH+cM5J05r
XJpbQMVPS6kGwUgH0SzBsKicjIQXtJYoMzzTuJHcNSVqS8oD121zBgusyGFWQy/P2ZQQ3lJ5Wllx
5aJTzSQwGQVXe7KvoW1210yyDWyd5aVEB5SihKiQH2k6FAGSxO4Kb3SM9CW1frAkwCajge9WUVui
zLyypNNhRErYKTeUzU8MatJG0MO37IyHzwsWWFg9HtiGpa3yz30onngPKXnlev+MdZpNp+4vd6Sf
0j5LylCT3Lf+jme3/kiaHrj3zIHJj2/RLFXUe5WnB3rCHq8GQR4J48tErg1iOjGpiqd+b2Ax149h
i3mV1/xcGAMim0N3KxRVKt3tY3p+xUFAjNKUWcTja3wLN/3e5hZxheN69RxTqi4Y+vmNA1StOnfj
GDj7whEc1+IipjIjWXoedelZ4OcNhtxXgEmBwHGt5ZnOwX0/gzTRFpLa39W+faphmjTcTP8pgejr
c9PTbggrviBS/prAi4RmxmJhesxKo3eAqP0OCBxW5NehzsGJrkX6j3p2HxNjaGntx86X4LBDFkqv
N7LCa2oklH+Q8F2FsggpvbTSd2lUi1qHvgS/GpgcRatRBmBi8aTb9YMhMZ9PPQ3J4IME42RVJXhB
p5kRDWaLUrDq2xasvJl1dxO3roegCi9l5oHhL89XNGNN2tPi5UE11dxGICrItcz3qDWYByOKazrI
jxmlr28JaVBanCOSftsQDn6yg2ICrO46PjpMHIMtrK5HxZ65S/FJ+cdSrv7DdnQfBmw5SpKpdfII
AymDW1e1juE+Nxdt3Sy4M8yc2RC4pxfCeuDhy9abWeZZmSZ4u1eO1dTDdXrvt5XUN54z9vyOi+Zq
1MNtsKS2jPw5J9fvufC34ggqBsKzACgPxjk4zD3fs0vuOM2SWNubXXggEAqjwdEuvcjizcMuPLnO
rr5+DirC2DY5xnXrfOHjB8XuysGQcePFyiNvM1a59T27f/r6TEUckYXEqgLRNyk8lHEUS+NSYpQl
i8mufIqCS8BNcU2iLmcuHMj2fqVeNqabV5G+PZXaOigyNizY/ehzYoUxczGqFtVgtFByzvc2BjKo
fOk22oJGqThpf15+RpFozTjTHnb0XjKhJOuqdmI55mzYx3OK+jNo+hO6oC/3ooOOaC1z1Ueh/uev
fgiq/onzRNCW/Fk7NLBuRrQH41x2rb4v6z5m85Gfhzo+t/q95Z0tqdKpPk2GeYUMlx53Oyv/fz7a
oG0uYOaCWetud7YCKs2HOvAYwM7PNLmshXmf54LrE0MM6Rrg1v5AnPITL8xVOsEOypPCRqyz00Nj
TP9XtO5iyLf2VbkAaqBOHaSGJTnFiDw99sZJ1dOZYB/BysiDK7kr8/2gm/NL4TVZAKBClL7C88+N
hifPkIei1ibqkyKbIAT5NgxCSW3CxSPCjDqyCvbR/JRQbTGyup6+gLcEaFAc7ab1PzfUUm2UEbFH
lHQl/JkM9Z16S9REuKbFQXG+3NGOMzKvB8IaC0b+h1R5yRlaQN6A+DxYICwYYKjJfCahgh4reGH3
mK8+B+35D7V4dmtoTYs+rL0aOWjDryQgIhX+tGXAGZWGjgWAxxI+MzRwRjoIvUopTIB1eIc3HLNm
8LWS5vJtMmcDJnIWfLxbCXJf9SLO2ZeZiwRMu1/m0/0HuRUhOZgV0GzEoB08QcMz2dvfHM8BrEMm
ymGiAFWwKKxR4Lp4DMC1dj5Hdb0bmI55Gi+jliqHcrHz1F4deSFYBnoN8kLGJLFQ0fT3Rkt1Y3s5
ZY2oXubEjrwmtfrFytTJ5iVBGrUsNDr7GZQOW11xONpXoywB8V99Ao2ddIwAgLVxq5x+BnvzbNWJ
kccZnFPdt1SPz/nBEmrFoP+Cq8tY767WrIdXsTDWOsyDz3Ei2iOxCgsd6i6ReB92cUaY9vGSanVF
iveKwWhFJ3r+td2AjfK4SATnAuE3iZHXnqClfovlgK3Sxly3Qpy9RokgD/FMFPUy/aS7O/iDvMsZ
I7mcSxrpSG8AzvU7PrE0hsUf8YT88N/W1gwMBhh0ZefDDg96oE/EQAKHg/ljAe5Cw96yq/sLNUvv
LWoI4xnZeaEp+LdJRXW0298ERdHTjRs9ID6SqOtwi2quyZII5VjEfS5d/27JqfIkdCNe/V8jxg+F
Q/IaeJch1joe2No3FebFhu1q6Eshjgx7kYrC6pM59I5oeqshPL6PdVs8C3HQWgalTY6cszTjSvap
qqVFs1FC5scUtf3sbA5TYsmEwlVs6DvF8sdaBCpGAB3z62V9UHbpWWNHcnevh8XLrKipV+I9/+IV
qBSAUhR84GEHW5AaAcmCsEMjUTxUt5AwcdiAhiTO1t7osS5ipqqNJaqETo4FHULgZTvou9+7nVQA
cDC7BZH3aKrXQtMe4otYFWNH6fkTjvCf2bUettPQGN+UrNjsiBW6S1CsJ8swAVB4mWMjxpxrT4yN
bep3jMTRKMxTZu2CEuzbp+8PcyKcUlLCBLlxHuYVYNgwexks/Pa27la7myyY1fSMheTNVKLwzO2N
g8xFOFJcC2YvkSHlOTTi/VXV4ovFCt75k2nqlK9mpw7poKlBBmzj5jrPB9qMxRpoMmm3pHFkuH3m
19EZ/iwNcxOJ75TjqRYhjvPN0tDuAVkODbDo+CQ3GMRAaBKIez8/brKXsu7PFxi3xF2b0luZlOBf
3uK13rUaHNghIL8lyikAj6atDnjz0SgW04VLPZhYn3JDJ1ky90SirMarZclNmnvYKvh+L78W/k9S
bTJMDZq7yvFBgbPEJIgSjAm0vwi9sk3yA+NVgjET92fu1mOcOdhQ1JGViQFvbmG0rgML14gt7Pm2
2W+raP3YVQ1JYs3vzpEPKFShOfuoQOYrFxXZTSK7Bg3EcWF0YMBgL3wgoA6k7lqBRP5Pfm5e/HTc
lu9H7OfMHZIF7sicknWTpoiVsSLC9Up01xmpjxqSvspev2tkRFj5LuUwzvJP3pMDWaDMt5AvUfkM
XMeft200fV8AIw0Ij9ewIOd/UjV9rKNszQSFEfED0m4+eyHz388/hmJCuJOc/7KNZafhKXr5a6MR
o/6FGa6wp5yYmyiSxmKKWLkGwzWmQWfFl++JxqL7+JW4K6FaG1U0eXZAtQxoCXmhaOv5x464uQPl
+/+M9ZsLqUL35UvzcoUBLmp6IUMB8fKc9e8FbFu7Ogs7/kjA8UDhUtW1DiKrahyyTvIBXfckK1M3
UgCZHAgoEGRdPspOHtaPLB8iI5EzmiiFiGrRiY0XtVPeoLmBgXI+noSOY040mepwdwKXJTB21qC3
twWSXS0zWkMyjQwLbmrmlDDNoqprfqftkOpv1o6Od4aaNH5WdxNcCVwYbkrJgK9t/2v/vnA+Aq8F
8TnEDgcYCzkmz+YcpZ20BjQexRbEGdQdXqWRP+R0TqR6XkUT2Cf0vmI1Y3zyXTnO9Wq2fPe1Y7vW
dTNqEQqymeFWhJw0ds1zf1UmzwJoFTX8EdQCEt2pMIh1ykgvbaQ9mSttf0iwZnKwApM6udlofGDB
0SQSofF0GtFrS8ZHtkNKpTniil2WMlEWQQ8NltM3RBGwlbcZW0Slvxq44/Thn5uOwDSomtQmUKcw
lTA5JbWhOmTZR/jn1IH/mz6x7exTtPLrG9d83gGR4nJz8DflVCSgvO+bBoIZb8xvFqbENjw9tyCR
fTZzx/zBQZDQ7NiFJrYvG+2gO3aCzesqnrVwh2zbkJ4St1Ay6gtUPcG9XZCTuTNUWSrOuPQLz+Ze
h5T4mqcOVHyArSf8M05NKROBDD8R/xkMC/Pvg6FKhRKfk8G8ZVArPM7n2PT5qH6MxRLSdhASBv+1
sz3k3tx+5MKiCEGjRxYUaNkRtMamumlrVH846Yydce723Td5inbSso8eQXYUwbS4tybU1iUQiwRG
9/1kA5rxOPGWLMTBCVhMXmZ8Emv6J8rbufyRG+Onzi+iXz3l07QjMJY1jH2EYuNj6he2jV1kI/cW
5IdaKMJBoEDNfl7pEEh0p/8SZvn/LN7HsCUZj5zBBp9xaY229+1DR0ggKI1Z9Zwafs6YM3OWuqJ8
ptr4e+oqvUz7H8bTNl4m1iPHY/MQZ5ehLL9C5/QgFaa+4ch2v7hDXBVcv0wpnWNmbeLpVTuEcGx1
kh22yUDn8hIyQYpm+emwFXg6F9o99jfP1TGSHyhYxWITfwDwGTfIREsvEM6g1V67B+3a8nj1q0S/
nJpcEqkxk0JF4rOTT67V4b5T/uSt4HF1xUD7A+AJ1y3wZQvB9bu9O1y0nfz0IJwEXxU4mH11Sibz
YdGcIZk1KEuyWQQSnO9f+xKrhbe0FMZPgX66C8R0L+q3J6tsloIies416Uy7zbHhvwqPsKKarvJL
qvewmoD+nGc3rYgJc8xunkLwqeTQUWsOGFk0uNRWfKfhH0mLSpzjB7giAa3W5+9CnlI8WR7fWr3x
ys5bVyD31yXAzQXFCc2KZqdZ9m59bZjqw4AxfFN0tGoTn0Ql5KeLy6H8dCUlvRmGLnyc8sw2AFQY
3B7suAAiEvHQuVy5UZ3ik3448u3k+2w1kqHq84owosT8qpoc4fsdXSDMyRyd+FvPOURhF3nZSfht
qAUI/DIF/k+m9+7ErCiBauFKxwqY6O1phHad+2zqyrtOn0xCnkpeG4FXPuQ+h/vAmHGRPmSN1sPy
zVuDavEaMvwtX/9h1jRxJBAMP9u9sI7id8K5rP49ICqUqNNoDUF0+RboVJqjwTPR0NaxnPkMdw2H
ECdbnF6io2qUcAOjxsyA5uDVPlywzGDhFK4qTevXsrPDy+KRn9zQsAjlk+pxdV7rjO84cdFNNlWt
cWU+QBmix6XjJfGK6O47QQKC0uxP6gW0cUfvvPiCvv5LmL7RC8vsCotvw9zmxd+rK344Y1rwhDD+
MXfz0GwTWYCZkNH3ww58agyc3Lng3hIfCHLTO/J7c9x01a0XXo8FGzZWkusBveH8fkCjowCA1arZ
Kz2Fo8sQbXZZU+/163ykJmZiT3+xC202zhE/T1PfR+/Jzs03dNvvEZk/TUn8IrLNh+6y0s5ApXlU
wbl2pydoHVG2ojTdKLD3GF3t+BtMJTWK42QyFTudMVcX82bXfJAS+StAKVKdYGJqiTmC8v2F6BF5
EC+YSTCnZrpfeQfzTANzvfnlGK+v+1xgW9nrTkOp/eQfo0g6avCdGuS9a/YzYVLoPPCJQJEi3e8e
1yWuGea68aawmfypnZ2/iDN3ssehNZtEl22eE6QvEuXiUjMBav6Kz/4nTu4TFh17mnTPn1YDTVz7
HO2hQcEoQS1VrDtcj5IuXq1VHDXOcAxitRhliIPXS7l1ZNIe0SIUcj93vjPnwU+3QLO67hiRgvIR
e5lULw+tlCid4xfgvTj54rg6an651YMIyGYg9oJ5hjquXIrLwdVgDiPnlTCrElivHneyZ8wr+9Nz
v7Q9cG0txXw/ohOgk1YHUvrYS1tqeOQak+ix8hYqbzHspyuM4YYu5hDSQWNr+3iJCcD231AfCDZf
+uYNz25gRAXvYyWNU7LlFxSX39CmojfdLKR1rCCjyfvRRjFFQyTgl5WVnhVjsRbMUlUM6WEt6yDJ
h6auMdjeuyqoJ/o03avDBkuubsCqMJ81RbfQ8uIVCwmbslPdpbbPVZVzR8sd75NVhSsRDn8Weisy
vI22DEKvFPK3HebDr9zQJhUn7UJRf2XmlmICpfr9ve0wgJwXrjTWZgfdbdKQoYQk8CSAGhFXkk4P
Ks1YAaShg9mRJY9oCkSC9SAhaGYPCrDc+ublR+6xFXIMfptNpWWEbaHys5aVX1TaVZq20A7yNtlu
KKD2DBEQuBz0RVQ0A55Yrd9GHZHrpqeoVClKzG9KyGD8OZ6bCyHTVl4hwy/W/+gHsbB6gWxmg03R
cU7JvvjK0u//Isgynv1WlIg6DIpliBTP+YQS61+nA5OJsBOUcmge8TQ3vNQ1kCTfBYoRkEdlWsWb
zjUJL+auHttq+XM2FmOCmVu7QFuXrvwkDuxVBUCRWiSklkG9sQWu5L+4rt4QJGt5ggPEg8eGKVdm
+EEm4NDH0Vy9YlcreHlrpPIlFLMYbSnPe8W8U2FIrAdE5l6Ty4mAbh7oqA7QDvqPq283Jn/z0f79
05YvoecdaJHvBzqjB6Ib2lB+BWFxMP1155jEXQoR9SKRp8Y0hK0rwiMRgDS2ugt7AilMQqhC+d2E
g2l2nTU+qHC2ysdfQycRgMt4MGqdspFTWjy7Za3KGi7QeVS8qPZ3e5T0tpMYGGs6cyplzFAh2Dxc
FXnOR6DckC3QitjHRk7A4hwPWffFCfX6Rh0cVA28/mw1L5uRwD17nto7yAyOd2pdIJfwvKf7nFAu
Lv9E0jpFYFhozo+ehza10IZlrdNGXBF8kDGH7GvFmF0kh9btRWxeneGmQR//PEhuwFL+xIrozNXX
xMNk6RRKUXMou/2jj89Pu59yuAWjIeubF7xm3adK8eLYAXYrjULxHcxGgW9QFfrVpass6oB8F0YR
t97ROnzVh+ONhR2+OFEhgp1ADyXOXdHXHRpRfc9Q7eaUxqg8Z+bLCXMFzUrN65n6vLeOqt9RhTil
6BDYq/TtYgrBO1A+tuGTRc2L3au2H7m8PRIG0qSGh1luyuJ9ucsErp4cUxwAFEh9gkQhke1GiF7W
gpEOT4wBSiUdv5f9d8zUlZmA0QAV6cLH+A3aV9ONUjKfqcbrumQx6EN30YhjxP5QHqnI9OQ7+REF
tKxzrg1/7E7RJpZ6acwjhKOrlDSh97Tgd5wwLcAcrzFtsZvxnG91xIqEKC+Lh2RGDHKgOpMfGeaI
izWrZO4/6XJ+cpgyJ9KX5UkLGabYKyCh+mRlYnaN2mCwpl2jsMSVe/22A9wDMLEsXF2PgPNLE7mE
52WvCcva+7pe1uujekm/Dh3XJod9bi1Vpy6NNlW27VmsRO2ZdvLcTzVCaUDJ8Z6JASfnweNBSJ65
1SDsT/2Xj5WsVDNO7qA2d2Wedlj7iQaCLnZ1Ym2ed4NhTHeX2wP3L0Br9x6gw45A/VyCxu577W3h
ivjK8HtUXFyCWEGozrDQVaOZvsonQjWoLXgdqs33iDR0SqoZUdtzNMSIaJ1EGkr2YdLS48mKl1bm
q3Rhw3b/zbAbfLExzTEonZiN6Z5razmEIIllNIxNc+RoaPAFe2Gpx3FDLY4D9GuP+AFbFskuCKBG
nRGbUhNIqRNqCJErTC6eKUIZ+x25ZN80luk11jEmTy0ZHgJD+F5wdOggN4gj1XkxS+qMs6+HwAk5
0nEu/UCueVbZglKTEDoV72q0Zgt4BMYSa8Sl8rYc4u0DFb40tlUkP4TmT8IGeWCJK6Kn6EiA3c1I
Aqt1JxbapNBqN2Y0q7F9nSpWJbqUnEQAde37eYq7Ze3ovOaQQ8sEDiC6gF6QEyXzxGsLbmY9Z0jk
VwFQd59YFwnN0kOkO6agP1DuelCkHq1Ox5NlY2qf2J9A4nqCrZf+MA5V76khaDP4lHJw6sclptko
horOWqanE8i+HqOX1KqJ4kgyBxay6jQFzBnLHLqDp7DEkRhyiYwO7ypY0r812yAhh05giqAME/cN
CAoeBePZ0ononaMHgxhiQYZZdcSdL6S/JjqnSfECoCDNnr2lrU5rsreJhmH6RcqME29mzWOE9wCv
H0JatmyjA1BWDfFW9GD3CwnS7sdg9OzJy1W3yOAC0c5R69yQBMJdSzGbffVha96oR+hLiE+9Kecg
ybBaA1khlOfUuRwNvrGu3SMq2GN67rgR+e7oY2j8wqmvgQzO99yjEwDNUWxZZtEU0KVJwhhKf6ep
4pi7b8fastOC4q6ihb9mYEcA2sVEJfU8+PXUzk1mDbBD3bIIznC/8LqH15gf+IK1tjjEaliYSfFN
mQSMBuHRvV9PGuv2lx9XjV1RGTVFbTT2BQF0a7bhCw8uwKyq/cdKhKJTEk8BtCuK9W0nCwcC6gXG
odmn4r59P3Vd4I264vgb9ByCkxsBph7f0sI8kR2z4U0BRrilPuAWKM3oxrBk2cazTHfDTfQjIlB1
k1qNcdsriUZJIOSmXUggycoOr8F9yeECFF/RtYPKPVSszDpMmrzctAuMW3fo/H7YKNEEjXJlR0p2
AhDrT8L3PlOYLt567Q+lKDUh79M/I3sLlN/bcoLqNCcVMU5u/y8FHV+lxEIS7EEM2txEP8639bpo
7nUIyycOHExwwH6DS5e+Y/B0h70unWsbNaXsvttM1p/4mWH20nPbL7OuZC3lyzoH86794xYZAgL4
V+k4oCrT5YWfWURcYj7E9PqZk1Ox9vAsEk7ma/DtFbLyzINlho2ppuDVoSSwiY+lcvBL9qGsjDV4
UCgr6uq36iW7rD8qzZR853JiLAyouO32r8n7V7wqtrje/ILEdjkWC23XanSjlViurs/ryPYz5QmV
jsnJgsM/QB2Ok5qV7Lq87+w2l7Gm11901rTPDZuwU0NF7oI85EIzeW+yYRoVVKac3A2O7AwQiGmQ
LmOTlQjKQeGcnzsJPTuWPslVpV4WRsiJyePsnUImlWAeyAIoe70ClP03J9LecHC1WVaCiDprMA5o
CCBEIaFRACZpqDFolWlbnkVsNUuZRijqXQ50OaWwzqbg7HdlUBNtjdb3yafZUpnc3vAywhkYCQ6y
Tz16Qn63g7HZKcoI5PHOr5xr20YRHnbingkK2pjseMfAmN6YYy2oVwr3MInNteL/gEfhmwlf0m6z
Il1xJeviSsCUu5R6uciQFUOAezy1BTsTiqsOFAM7u/f71yRy/uq/kyz1XbJQgx3w4I9V+aegXzot
kWeQ8doaWx/43aVVUZFpVR1FSlrHm9ezvR881sfQ8Zc2MxYwAdzTwcnXaR7Arpw9ZGOEli/8A4Vd
bZoBO1VIR7JZoDRjj21j6aI87iBO0Ov5AnYoCFs6EECgz7/oAaKwia231PBkluJO/82MPjvvgS/k
yW0TzhFnKZPccA0YSlrIGO7BbWVkRKxQwBrbYJnj/wluVGrzp34lVuCZjvRStM/GMOcbjiWacPxz
LlNplKoygTPha9E4sUEHJRJvHF04X60YFbwYcLFtYbDBuz/4RoPmqisof639qYGG3PMRDVblHmtX
npQHglfROYiwp+QmIBFlV1Ze6zi1+VaApeOEXxJnAqcK5hAMLoMrfRcE6DEnEFGWEmNmrzLc75j4
Vk2hPW7OzO7aInkvEtqTIGz5udClVh5VSZ+cMdtmRvtncST6CZ3w80Nht2pO2HG2E5xjZt4eovgY
rUVcFN2+k9w538zezY828T/AoLTfef9PnWdZABCK13gvzQntHwWTHdKG48oRTL2efOVRFe9tgWF0
mHVjvVk70zhCnvWHfyg9vi02YOkbu1X4L+MmO8trno7heQ2SXGdXaZ+8gL6qebGZl3L1WjKrBGx9
G1n0u7+BkDd+64L3Y+tzIu/y+TQLoyYvIFiZDqamtJlk7fErTfEd74uQHaDhw4v5fWedFFqyi/QV
ctIS47NZzK/WSCGo+W9mnqnE99RCPocmZKokwtRldlkeZJrXgYGtlDLfSeyq+M2SFiF0W/nzp676
hFkO9G4b9ie5OnfG842rgvJvAbg7hPLrma9IylK1Vtx2aSu7W5T6IkTyN4IBCKJCDjJqSxa/Eq97
srUA3dFTVFGTplVWi6QxiKyP51GEJ3jvKfu8BKJJ0y7PK5WxLNBPeYUg5pL1LqZD/iMOMQFV/DNR
L7TH/00cJRrsLB3eJL+8afW4sSV6p0+V5iwujO8T9BMvpp/1tYM2/uUpBmHGaUhaR1O8aFqxp935
xdpFHdzPXUIKG5mb9LegDNwxqr+kr4CXD27f4o2KSk2y+u2RgDHQEqPLRbYr0Fb1n+w93o5/GBL+
cvYZrzGh1khT9LMo3q/1yVnxRR762hFOd8A/BmaITHqM2n4PhTrCPnUFpA0gzxGpM+6d4XLW45B7
j3iGThRIpNKR6zPgaDK1g72CWn8ZC/8+9RqGxPxgVxByZeXtBHkZnulZbpZWoQT/gpE7q2pgAgKM
JExlQ7Ycf7O4L4R9oiYaahcT6dAZaVKKAN+fpDcu4sQemlVqen6NupiodCZvfk5Fbz7bi1Na4Zno
n9AcKg+hqmIGf2OgSNgqs+X8Od6ARkaNjMfv+710shGiQXGe6OGblENnvmhXJRtY2vzhts7WFC5M
lWx+sY5eijAteyKMIT9iaDh0YH2XG3AbpsqRcaoFAAXofzbRWtlwU+x7nRPjElemtZ4LKUB+ib+j
cad9WJJiCIZW0d5gs93KfUe+NBgl4HLSVGLa5ljj/M2GmhPn+dvSyZznRt7Yqpv2qJgOyLXyKeVG
AyfDZRw5N0f2tEF1f2EDwWgeUVFRFlUveYxdSAhM9kAAfPNbwqbt6rAblZWttkXxFg5y58lcwHy1
4Sp9pUZBVKfd5h8xFuovM7pc3pfhK28qrSGi/6mKMvAa2CD7WxwJBG7HdMg6+pILfdhiqX6EtqiI
Pj7ZOetrGCqgDb1xwXQxim8jfsWRRdTrfGKVZAvjDIPbS0pYTp/ZfaYkkW+wUdckdnPaJZTb5xDh
amy72f1ovc/gkhH5WD2HyrrabnrH+99PT44ZxucNORzj18iAe/XFn+qbVzsBagUMZcVqXNUm+TZY
x/cuYKGf74pk+7XDkqC2eitWCTxsq7WWEU2BOt0xu5YWa8Nbvx2qu+JzJ31eoQGlk51mSy/N5u/V
12UVIt42nGgCuYjqMU3ks75wr5d9XVLuOoraElehpPzoJS52pMAqDwIXSN/ZRPxgEZ3E0234HWN7
dtdzOCuaCRNVsaWHuW9BbdPacEv6sq5EPXKO6GYdx0HdKolLW5AEybrcqr7xe9uSLZ2zuCGUoCex
/CvVXBF5jPlHGorEzza36CPkRc1fFhUOCLA5IXYBnP18hkJbTlR5oVlehcewQ1wzLEMJjbHt1piJ
UXfZpZ1fTIEwCBGiMNdvdC4ro2b6yCkbBHM5sCNYZ9gjo8d+6aK5f3VmwCgbyGYFsB4ln/q8aJVr
piRi+vwlt10dk6hL06Ao4saxBVVgzpop9TvONsYwX7uAMJYWL8sAlZW0G92JBxc5oiOyBdR+fheD
vec0KTIDkJqFWEXgqkwjKJKpRnxuVLIgXTawNoVKqXZc4nKB3YMDpI/CwVzdgim5CvEIQXJ2wFrC
C/lliXaMFlXZuJZqqoUlaiK+j0J3aQZZDNwHf+ldcdJ8PYuzp6tvr4L1ftNo/m8TwFDYwlrfNZ9r
GDrEzmBksA4JNUj/yM5MrWdWZ4jbJD/PJGSER0IRyWWejdsGiABrwgfhuwzlt4k0nDMWoQuCPcd0
xHHJDxQGkGDRRriypp2niVrGesQnaTVVZhZzxuySkudQr4brAvUNllsKXddTQ85hg6ldPt1XHM0d
4Plrg3y9MFfB275uVHdQxeYPJTqpnEnt2lirEAfvXEt8voI8uEojfNrIrh29+v5467nZW7GwXhXz
fsdYQT/lGy3d326Pu7NO4A/0P0bka0VnfncDw0gPxKfCYrhegG/qRYlzxCyYNmAFovYSRNJRWUvt
L2nOH7C2vvlCTGPl2kjHYC+APXbxJlSNMrYpvrEZsiR7LHxcPuViaZJpOPctRcju2oXk7DWbmibP
Lf5r+t3cbnyFfLXbgoxRczU/M1D/zPjzpvlcTfCJflxngDT0wkbsIh9IoDxux90AV29C8wpTcF0/
RiiDan/Q9HL0tcmrydHSfJI61sCZIv8Q0ysFzJKrUTPtn/zZQ/6m4r1kYW4nUCQhK3GPw7X9eRSX
JR+EOyFGwBktPEP12Fx2jrw5Iv1Jr1MDcql3CkZMRdg/iWY7bzc446BXMq94WrABrMnXA4sAR++k
3n3qKHlqDZZu70TLo/J6uoGPI4VaCdAJuEZWgChSRJ/r4b7JrC1Kw7UqMlc4Aj81ZsE1IFG1SUOV
tod6tiOHj+qZLOA/OOtmGDmj9R3YqnuVUd8UMtN7rPdO8rj1MJVWL9gC/Z3SpdXzJxn/8r3znVJg
rHwF9xUTrlff3X6ir1RkIChNHGK+YhCbGZn+JRXHInGVWdyFb39kCVfZJpliSl9KzQxjY/UgyFO4
gYdz4xtKIZOBxZ6IcVSDgJ7n5bcspzYrM8JzhIWDxzTaWr9bFhp/ld4AHSlgBI8pIYLwmouL0TA4
GV+xYZx01RA3oP20RaKvZ/eTCs43GQ7N/EZntd58ob9zAnI+DxzVsztxKL6gfG9N5fa8wH0Ud9Z8
O/k24RVeu9Xc7oJdrlnO2irxpHzeMZoUMCZCkE2P4usfQ9hrxxtzow8ZXPIsq/Y8z4K5d5Fixzxl
60+/2n4Hn3lgB1EiDRr+pVhVJYBTpK7qqyzzQ/ZeD9V2/ykLAmTMUSUE9W+6C4aD8vGyKKUfhLaH
zceoT+pLs7+B+PSJGxErfIXOJlUPhriU/6G6fLat8iljihu8kBcwBH4EFcc0IUIrJQ5AhWlkWGhW
7qGjrytdD+GI4SdZqqNl+THSAKu+NsVIYrHtrK3jfilzBnIWoDvbwjZYbYnhn/ZEzcW0doH8GCbq
mXsieB0WGSyFBfnFeAg+m0GtwlhQMRuyBQnO1WkQO6wT+JcSFC2uJQSbvEzs/bDiSbXRF4GPUEyC
O0wO1DcZTEZVEm9Sc/cvm7NE1ALUnKD4A3Gp4ijQykQXAe5s29R348SWCvkywfFvbjoCvDsI7s7z
9daWQFjAGdLVhrfrGwmcqSfPDeB5RwfKrCX8fU0LXy/BPn0Ko1XsTsDc8p1oaejCNvCLtwRiRwdk
rLVzhcEefp044sQsywOCK6bk7bVTuy8HFW43+xMETS6NQshmrnn1xRfhkJZuMidt3TIDRx7u6BvE
dezaHWc+kGCL7WoLdnxDmeNSrcN7plXtD1q2SCA5ayv66+5RFcUIzsTZM18iyWls0My1oDiVU3I+
t1vm7OS2XJ3+whc+lerTUFUIe4TbhsXPAXsV8IaPeEi0eRUQbSjJttcNzyps6I6YOjazJxu5a5JI
vHMT5UK8HBMDUHW49HjU0XhYM+qJ7t3H/QBOokIA0Vgdy7lxPpV1ZA+vBq3MB01X8aLVRCBRL713
p20ByBX50ijIAQa4yZ0n5k9sDOuJ4YJCXPHD2y+MWpQlSOuTPtMdG9q4WGq8UO9Rfw9IaTth6xA8
so9cu06RPl/ZfSrBkB5z/VRcMDnhinm46FD2rTU4XzHGplqcJR0TpZ0EOogAI/ChqFtbhnbntX62
PqZzh8Lu4Krg+lXYoOwfTvBhxPOv5Rc3/8AhYluGYwiARrp8M/ZiTR6wfxtvonk21OT/kBHuQfNl
i9w/kzJcZ9S3FykU4x7Q/iXeXqIP/cpnEW9EJgLQvQ/xNFwBTUoqVvFtx/xukQLY/usZq8XeXrwj
ENIaZvj+qw7ZpK7vtf//0S7G3zHsmv4frNwiXYy8n4uxyuwsSzUTJNUwX0MEgeJb3LKjqhD73sEe
4o3HLzvbWUQvY7jWqjEjWXaGpPxPvfM5aKopnEQ4SCeHLJs6pVRkLOKJDhvkyFwN1huuzr0EM7MA
nBDExDEfIGUAw5Ed/ONV6ystAfI2ZVkGKLYkupxdqSBoIzPlKXMe+owlLUwT+St3XIYplZhPkQSR
6yMzD8VOiZzNCqroE0aWcIdNGF7AhSgXzZjsuDXuJRO0hkLDpLjKM3Z70ewuTZBtlX71lwSCjGEB
RlZsvYgac9Rzw+bjBan6SOtK/Vivj7GH3YgFVBb8Ivn9YtvKPHf573ZQMmgFrreeBYZf13hZHv1k
rSHPazGUdyqeYPpL65DL1H/B+VNBPjPY2F2RK32tgt/p9pdiGnOWlMS8mAUaenM7Dx6zQLmEOCTh
HdqBT0GFM2doHGGi5ex0XdMlYbkZ+SvNrNX47xpzRF5LwFSy3FHzWhhWBPHKw0ZE27dOaSzkY9DZ
H7GV3D17r6ZP6xDbcGoY1MjiByUcOMZK5F0hxoT5TI7OWfQfMEz+3XkXCazNtuDoLyH0O4hPkP5C
jtfaR7fHVxvyZZhNJNqWWVAaK+iMr8Mxxutl29xq8OjIm/FqQ/TaNWsNqzb91j0D7M+ltIxGQMbc
viSbTJdFrcDht1GDsZ9vsrZS8T/D/LXFocjBsf1fm2+keBqpLkL49sUjrj88/kyhRACx5XgY0aIS
x8otboZrQc+ZbYJncGhHFVCxsAGnf0BZCqXBwtd+WtVVrPb+Gm50yme5zvgqq6KN7vIW0Oz4RBsI
NnSezpnAb8Kvw3kpThvYHa3r6GnAYO9zimVW5p/UCPDdENc1XmXhp/QjvXV3VF/9N3+iovzGNaYM
/tHg6tc656isyj0zxFXqWlD00g34rvv3+YNnaeCjxx4K44eO1QAzjBA0/l0xVpxNfcMQJMy3kiNW
S35+Wi+5WqEqGcSd1D+BJqzxhn+yUasFrFij+aDBWtRpcOAPzYSgq/H0la8zt7a4w7TNeY9x++Oo
OMtmq7ygMQLyEAdlentl9udSxnUzuCnc3iQMkaBezZCbUwAhVVpMLEt3I3z9qeySrsObUJw6nbV5
u53i7ZBV/bUH8fdfSsndZw7b7o04vLz9qqr/tFzx6Aa4dLlwYmMcoh6ck42nIJGFPNI6LLA8DE0t
0eQN9n6iSrO534HqmhQvtH/Q4n+4fWbj5AorhIr1TsdAI556ot6NLdjK/rR3m7umRDEnIUMxfDLd
yzkTVWvucdVSjMkykzYjntRKaXPrMBDpshvj0H3jLBzEvMcbk8x0+zobsKU3C9Lj/7jMKkP+qvoN
lg0DVBmJkEzlO1B6yxsWD7dzFCC5C+gEkYHo6rhZ6JlGVgqcyUajvd4mvesHtgSmIqF3JQDQ9yDn
yIvCItPlE/bexy+lyOz/Aq0NkLdq3Ib7DIPUA2IQuXQ99yBbYp99E3rEu1SqIvGzSg098khHzpiA
rxnYqErzZUOxuLizk0HWKMW16ljwDdtiTghLPyMuYsOIdVBJ2cV77vj+veu8nf6sjDo5Ki1E2f0R
w5VK9atQdmIyTGIqQVtSn+cDS3+5qFh0QanLCG2hEsQFFO3xoKT1Y+TCIyWPOYjfBMTxXcu2hqkh
P6CBKwQqTl9QwMUV8H9xXGBwTPaAyFJB/BkZosdcVKNytTLKCzPVU0bfsjkS8Ip5hDFhPmiHb5I9
mIncyRXZUvkGcGiWq6VKlQHdD23S3V/25zGRpWUngnQyYAhhfdI8fVlXbhdz0ZkYMvSROpU0XF4L
LDopsPm2FqEd5bp00BGNWHJphppWxihf/LrKx/Espt0idBvZf0Uy5edgZGmIkPRwV6Z5f75/AlXX
rLfYJ0QaFUFT+wAWw5E2ef1Ero7hAHyL1ud4kuC11+WBUGXy+IFLaTbQLKGRLfXyn2ltHMiR0rwk
4u6Fecjg/snAfjZtV/feOEBc/OKanprNQUGsgRCIWGpkXaOjRy6KJrf3hpA/sklLgKqeDRWprF6E
cXXnqaOtQnDhyZXC5J4oEGKxxAOceG0dz30kIX0jNOPWwJQ+FCr83WRSmDzSS66QgKakgnpBFonh
7p7fb/BQisU/CBX39sDt/lWfMJ0BC0OcvrXj4d/UhrKtIstCUnCBHWitqE2WnnFk3WS01Jjj3hpp
PsN5mO9xZA8EQBuIDX5bXhl2jMthrb9Adva4t82zOarAuTVVnNc61oO4Uw/uVrae7xmkojZnl7ed
oDk0hEEFjM7PyMwdsOcCD8IFfjFf5zzq2SKE8+AOuPwqL06RjDbkWP4VNWwX+gS64NmFhwGCq6Du
NpCDYFaO8Dq84JJW7P8JG6MrALaXX1X4JkWMVR48l3vQH/SZYaSxhV/UO7o8RbXd2vDHYXYAl9rV
9q6CZLuMii4T9YDznQe5ZlZMRuM/cHjnzTqYguO0CFls32zuXpj5FpSMvRPi2tFQdfuUVGgRO3br
7Il3l5GW9Rcx6FpvYXezpCAm6C8jr/IYlwviG6MYvQZfyIh/eKlZcdutEKihdwWveQDOLsRD1FtJ
fng723g8cmkKBr3xwaaVm89DW6+rs7VeSibdSicHsHLh+ppLoxHYEWUBdKWeMBcdeCNf2C5QISng
Wj9ENMVl57S4f886ShTIq2+HGiXYNResS2GIJol4ZHNj2/WEsRZOsXVFaGEFgKszb8OmW2AJ+kHG
ucV5ZOodRPhaE0t4z9OLtqTLLqxG9AEfUjiUgL7Z5xIUfgv1pNBtDuepod/CildChygj8SShYntM
KiVTatP1Q3XOxlFg2EGzzo6kqSfqeGVN2rZCRoJNQX49aNMf+emdxK6k+LxZ0aGYPHpd0hznD532
nQPVHwW2pjGBcFVTNE9l0gxR3UGr26FjjRBIJWQpcWrYMDvaMuIcvWoLPjG0Jrw7aYOwI5ay9Meb
nurZZH0ErCRsOBeqR4rLB85gzd66KdzuFyOJBuG9WyXxmSzfQYEEHubvt3ZXG8pJx1I5T3zcj/4/
2G8wrcLMGfi5oD4QpaJ8z9DYcP6y/DCaYgEMaTuWqmVvtSsOFySUr0iZmb4uM0MTjwLJee3yV/Hb
gCriIFFp0YduPRLnEenPUbUgoWMh7TN8V3ouX/NJQuMUEgvTcmlg9uILKCENxTVpfKONuujw4vcH
Fev10Rcb1OGttewL9hvM75PEMgum7wkCcVYAzjXMOS25iBgt3mtdeyzAuEZRWAbAAc6RUGIq/bqT
ylVdur0KnG4Rk8Vr4H2Hv8bOZOJDllTA2Iz6oyR3W+Rql7BH5gkBslnQZ36fH9MtOXdWUmeySOwd
aBj3AxhFJlPyjSqR06Mg1gWsDEZWx/pNDA8wbIC9VJB9R/cwSapem2vOo9Ybbb7qNOPM4pn50O5R
h1teE+L/0WWEyjJ0sCmwAv94vfQDSw+iZT052hfqUJmCc0YeMOTgL9kiji9Skk13HzGGsMJiYUbU
68I0l1V+1DbhfzTNCmjOK0CquopP66P9a3Mpf79ylm/6ZmZwuF/NoNQONkQ6EqMbOAkmR28te1An
oeunv1LIOUbQjSB2TTWybDbQPl8VGMehh+bk9+meXr/uUWIdixRn30+ENoFiHepy7B+qTCqvLlMS
+CcyPV7R8xJ/8e7CmkaF3pJ8LLACv/Nl38zfbVGgZ1k4PTQScr6F8Yp67/4j+Hy9yWMQI4MGT/gO
to7RI7K2kWbFKvTpttROhIZyLZ0ugQMmWZoaz9cDFgYhpzxBiv+c8856T0vA/PxEJBtQVQR4K6oD
nGDwtxuPkCyTYQ0g+dlNKWqNECLyNGDZN+dMJ0axD92Ow0+jtUMXgDxHOfhk5VFCC/tvpH/G/efl
yawzuH6nADpuTQR0VrFLirnOfH1fyfedbHQ9fdf4HtNW3CbOYT32Uo5BYZc8X3D33ElFVlh4mQ53
KDiq1XGRVStyB1vfcIsQpDOzG0w656CIvVyV5yAn0vupd/q7ec5RhPjIufmpM54epdAaQPP1/YFW
hsDiBR5NjnlGLDg9VJ1UxDBdNh7wvymbcQbZRu7Vqncg4VgNP89UutTpkbpthkGbx+TncrNGv41p
ZDZNqYzmiOvuseOQYR0n2YHerLL6a4r+HSQVPENnK7bSu2vp6UlEvwuSMXPocslAYvB++FecJbsf
2bFnu2xCXInU9auxrbtULTCwIPj/MdINy7HCjdYM/CyzOFl4fBY373gOkPhY5HwXgmIpjjrZS06H
4tGWhXtjZrXXz/O5lsI3BCYvE+Kynod7Bev6Bkmoq5/aUpmWPG/dqtt+RGA23cVBLncGofFNcJgL
4FJCahHuLIe99F/z8OO5oAM6eFPUAlZPgIIcbfmC/HW3gMOMXaDAyFPQsKqAaaqp0K7oaFjAEKra
cMtdGc1nmghkHS0zmZLyrLjZBKaRgQOaGKrtO2QDb0zwgdoyzlEVt8UIt7D/Ie66tGX95YiCgqcx
1Y1KLuGiLdYf5ok/HmMNQHxq2MGHl6kk44+tPQlmrHFd5WLSjmZtHovdzz3afrOqLNj8Lw6YA5hJ
RBYgkLq8is0u39pi7Wpynfq4lb5VOwo2JXg3qY2w9P6AuJ+f2U+qD9p4BX8zijCkm67VD0v2upx2
GlFGBdgJbSSCt4JPCkCbJVAWvoZDe9igzP3+eq1XBXg/mAzIZnaeKOGjs85dSw+fmmlFPJTLpUE9
tpmjpaXLrjjSd2RYBrOY1aP/2rU08FOcHwYsy2iujmYBhISAF5dszPqd0oWrjMrboca9pMhVo2+E
zhdfm2SVfC/RXCq1ZaC+fcos5fhkvShc2SGT/el9/TomIYl7Y/p0UaH+xeUpGyYPjlnynQt2b2FH
kMqnLFeMFwZXKlft/9VK0tf9jstFhG1VzlbUtc1KgZxFInlfkAG28SpNSPhvN1s0AT/uqpMqZBdA
Qha2zlgC7wZ45EkXoa1R8oIVuJwhT/3U6WMGCiJrSMV9D7DVPKEhSH3Jcbw+EmjIfU8VJGF2QtT0
+8QHPLuuYGlS+7v9yzRZgKVHpGfGe05RlJg8MKXB3LN/JJNMBLZNAxSbH/J6F9i+Z9vVQfog/dDu
InsVFffYVGDR5heQ6VIuwducYr/Nb7+Oweq3fLKOM7DXMnhJ88i/b1sQQ7pkKI4CsUKCFzx+L5rl
lN0Y2QbkAU3yG8Zw6D17bGCt7PFHPWckOTrNDGyKo2BohY6iDaGJO2KsXxTw9caxA4cQrEgIrYJj
oLuEFjBdMzkXO4XOznmLv2x+UQrsf2oW40hqFWTGDzf3/VhxndTmAOtnJgu3rtL1CYujla9RQ3PX
5prZKWq9qtV7TjcXqST7N5AQOyenSHAXVpB2uVBcsgYdxeSelDfoBtMf7vvO+vUd6vWvNHGv7d9v
lWY/hHE9B6CZk9eqMXC7qUCbHGVj+NAAL7LiNFHT+byjrTUzBELVH4B4ZT8SF6yXAm671gyalnqC
IsA0giYaPB2MD8hlTH0LO2Lt9/8LlGE6EQf6bDcV2GBMuU1GnejDrERij4aZvnlnqP1W8SLeIPxA
b8N9U7FsRaeMoqTNPzbom9VuWcaGnbFsiGXzBUdRnT05gnMoKay0hQIaZMIn/Em6AsjIRvtOI6K1
vKGD/PAWe3htBRFPYxCaruVHY/bTkyNyslVBkNCbjzNY/nIc6mxj7PaAXYc/X8KCQQQICdX+dz7X
Tl2pgiZBPf8xavNLEv7GUqF69qzFVHl8ocSL6ZiBem8Pq7Tqzg70uayBVv4l9mCDTeH8GDCjq9HR
FPj2QDVV9s8tD8fRe4buV4YxYNv2LGE07/9K+rJCk0KxmACr1piUKHA6ID+3fIaZqeRzbnMScGC4
HusA+X53ABDXLveJgVxU3iyhnlmCFmZuqwFlkfdlR+aBwpOgnQTfp9znJ6Hf8rbgz5QRh1o/uJwE
N67MBSsJV23JrG087CNCD2bm4ndEAFLI9LyUyu9rdIl/jdF1qINTbzCVdMKc6XZftRjB2JeZxY4z
JYh6NutHhzEOjEGW/AOwLlLFFLwxvyeGdam5lttfJhMr6Li/TQHX4Ue8r3k1lswcqsRHkebWa2VF
RKiUZEyHQiYHvH36pssC+R2HbRzzIruci2PynLuSSARhBrSUVFYQRAWHPoIn/Q7YzJlIlsMlwJ2D
euDJ3/D4hOtkyqAh0KxilH85BmlBCdmyjQ0zDGLeqE2iJylP1Dn4vvND/SllKF4iuvu5EPCCtGU6
tns7O7RBBRQcKH2fdV+iRnSc8dB7mzXvD9sHLERzMid7GMIodL+czl3hkQonWhWa9JSxqNF7IESA
amnMGw/bk4Qled0U5JaHtcEtANgRcjhvOr+SGMuwpUcYrlQJ8bvKQ4WXXdBNjI5VyUB0o8PcH90/
saxFB1FuOsGCKLtnZGV7F/N+eq6HYt0xwalxrYoUHY+csaLfsq7zR+gHZLgWRPjKw1FO+2QL+7cA
EZIUGaEuYWN0UjsdWkAfi4UMBBy5nwhaqQ/utiTiRQ6mEWpvVcPzIW2J7zYxQmnd729vB76Hwt8x
FpNzQlCNbfB+gJZa7ZC/QmB05GVL/e07uGJPH8SpFqiAb366662t8FECwRfbJyAk26Ya5LYW6y0s
pL5GXVhjM98JKxPJ/NF2MdWadJLAH6kCD/5IB7q19iD9pGOFyxCLtrwvtKgDDHE69civWixc597m
9jwiPxpG/mJcOe+lrxlY6r52zp9+5GraKj4E9z9vFvBxaCjBJ8KipWlibz4xxO5AhLz9OsPkKyxM
JnH+P4rVf1YoZtTcpCB4H34/fc+dWrj8BEsB7LESgTK2kJbr3tOz9TzQf0FweLiuGMpbWuoHGwhq
3rA2bWVid7oI+CA4MvIWdYOlN4lOYrvzC4n4w6GO4q0ZTwfkKnfnugMoHwZsWP65pFIIhZtYzhuu
fGZ87IY922Vy7KeBGko8CORneXbVU+gQfEHUIs6QLdQL9gSS6jEB7LlS6zDJ2cYcKcPIanHbEh1U
mVf/f7DN7DrzYy7LyURqhEI44tj33bRZvFcdUInAFdq5BB1j7k1U8XIZSJ79KICT+esYYUTxCHdO
+X8ELgfZdNoQP/25sy5resCw/2ZDP9sV9/2eP4q9kefiNbghCIsWqXoRqk3L/xZbSq29U/jDD8w3
RjvLMnYqJZrcsozCIhCNf9xRvQzEV5PiUz6x0/XNfoHuwpDFHNdW5H8stSqSLXDX46C9D3l0K55P
q3VMRjdkSIriSxvaTHNxHUMBrxqt+sqTcrTNN9FPpVQLBLn4HU+w5NzmWep8jfN7YEyNHRf+bn3l
jPlFiTBOgTqMm93jAHQlHm8UyKmSG6B/IPfxTI0dEyNeeNiL/UAwmvRJ1yCFKOGdjtfM6B/c27Hq
ZHKklB/DBX4jlHgOksE5B3j5K+R23Eys3Ip+0sI8cyYazqsMEBt0YtPh4YS4hl24WEsFxHwFDMw/
px3mAao/+F2KRVvZ7M1+gr3+dToGhEdx8Bdw0RuboW4pt5iR+B6u7lKpP6ZCMU6FF6e2blozmEM/
hwNijdX2+6fFGxS9BKZtd7y7MRrSJR5Tm0hoJ6Mw5AIjOp34MMUPzKymZtFWWw7FOfngOLecQtRr
Wp6oLhJVtERpdBIhDR+TdLY0Sk9D5gtMvk6FGW0QszlFrH0BLxJFCsQC8PuxYHwAxssI9ajzhG6j
MXpuNmK+GKgU5RV2TqlWQIfEXX7Oh4gadHoP1WTEuUUMLsZLOwcAu2jLKYJAAHP2RJ0HyHjadMDs
tB0EtoQrWmfhxEzUVJMHxJgU9inLZ3d8xlN1qpzk758Ch8n3ZuoVF6Pxi3Retq7iPNDv83/6SpuN
mNs/qh5vWCAd0uRjf4vjzTgY9yt+/r4y9tvDEok/uuzMa8dbVf57g021jf0Pvo0CT+WO+PutP1xg
aAnxUgGwwURGyRgmwNrB87O3Nq1p0Id2imnUyMrr51Vd8uZlcUJGAginL35/b26uuJAb9aDGCXCL
VnXUemoJf6LSO0O2GwNHqlVIuEHDtH3xA27DHeABtokmMZ5nb7OGUxbJon9k1ue6jWZOc/F2OV+B
IkBdpTdiN1mjKXowL0c01EDmuiO/9/hBZFH9HeW0yk4y8HHZ4gRv/EQ8KRCUT/A9BvrKHZqq1Cws
3PvLcizakthWqF0I3F96i3P9dPq9Ua6KYNmX7I0OYRF11vE4zAwJYOhD1ojbiHjSdx/pi3kdSu0t
OKLmQ/GjT4IRqz0cMmoYBfOh9Ud4+CkU7aePeIZ7fg+aRRWrW2lLQrQOUEMSdx6MCQo3Gc4sQLVM
ilWDxfcAyfd1mNQ2eGAvYas8EWnY72SsRpxo5jU6dPKZItJ2mL434882c1OGGk8rIaTWSyiT8/qB
WQWU3KzTgB3kFSszfzTV3s/q8jAjFFV2+wWSt0bv1KFH8uK1wBOuFHBrsj84SXJWciKLTB/iqkjH
7O99AlY16GjSoXdsAKOURl5mmfASg/NWVco/oMs9/jgQjJeo6fEEHXesfSMcF9Pv4TteAdb5Na+u
VeH/1EpUWht5pACBpHPIVNuc2mg8wT+nkXfi2alr86pFeCI37MaAU6n3UyvGPUAk7X7J1uDKSfCY
DcscRVRZwL1ZNPshH/GZWHvtnjI0Q2YnhPZdDDPB/yltjgzTQaUSTqCs8wt7oSRc+hAXUap4BIvo
Qks1V3fAvvCBK8MExr6Mly0I3rNIWeuk51xnBR6GXYGAcN4kERK3A9cat1us+Japyie6aT+p+Fa8
rCViTALZ47aUdff4pcLUVNHo5iUM7Fg3pmNbMiRwu5Wa4ZxaTM7tUfUfBYX1m8ojqh8R26lVF3aH
aXFnWu5QiO0uwKEmzaHt+iw92QAImnlDcyYZDl7E2+ZZDPAxzGxwDlTC7vMMNKPysBjv/xa0ShF6
n2tZc44l0/fNYl8H3pB8OpZAwpQlkJUsQ+T0iJyxB9Uhu/GYLhtWE2/Q4+LOBVag146bV8D1JXRj
IiIuvCGJytYyax8CG40MxDfYloaR0f0B92kIAMOxq0fyCtYoF46lW/zY4A8j9TxsiL1fGgHIOO3i
2UXlmbO0nrrU8wWJNLvh7dNwR2YQ3nRrCw332G6SxytUZiv20316GMQQdcngq6SiJzz8EvJD9CmP
3k0jkMpOALPcw2evnFQfZ+oJCrE932L7LJRBap0bzqWSkbnLLuP8k0Nf+JpnFYrut2VyYR5+wqDI
SE3xss2nZQwzTlUXnTI913J5zOPYQeVpCrUHujwGvayAbHNhSw05ASk6ixnq7qvHlAwrzPHxAteX
JELNFVtWQCtOX4U1aS6/hwGSD7pSEC4AWVdKOWC5vB9RPma1gtGUbXq+t9oLM4Is9FFn7G7HH4iG
gMuFwZxmjGaxkdhny2HB67rX2hjFYEtidrPQCYY5vJ0vJD8qQgWGLpuig2M/XK1nXdUvgeH6zk4b
hQMuwdZFUtZYI4akvM/0fOxEiv8cNIRVMWhptyGo2aXdF5A0bVezr3IbCmv9m28M95IdhTnkAveZ
HskHgxP68tezlwa37kmFvYI78tuDytmfyqsKvY9GuoVEUkZGuHkqo+sxCKexIyKiKlB3gfFYFjXE
eM/oq+/gvcPrVpBmdIT3dvZ9Xa15BBUWmiN+8SBoAeS3Xl3ZxUc1Xm3H0LNn3i52SGWpobB49K43
fmGOFdZ+EUOpgVtgp5pRTi0MIQSygBcQe84ansOhzsO9ccokQWMQIYFwDyqdFXLurrzLu38Ib9Fa
GByoyplV2PyPCpG24Kt+1Z5lKnz8df29gB9NN80/s/NnuWLBaAeVVraGWqi4p/6uCjmGX7odB+MG
3LxRNS+4Uc6/+uuk0B+SbRxfy/nfzgFoxi2KJ3E/U64aHcl0kpJsvJ3k51IJctlyzLDCoGG7tsg5
nB7EEFkx6VLJfiUuClB8dUqNCr1szWZGD16YaVeuBo+RSEEUpiJGe/hSq2mAYAFgvNN5QEHdYTYO
Wmk9GHmawVDW9IXZMZakyzzLfQm9vRoEYEtWdKgs+nBhVMun1dV41eUv28w1R1YiA0lhdd/X/re5
Wu53pCapqEWVGBGzHL77fly2XCQsPEyM/zEOUb+NmbgmIsJxFSxctj/rB2JcI4twwoMttjJ98X6t
r+jD1A27WXro22jBvsBgUq7M1l270Yn3Ou7WiY4D8jYfQo5SQteIeKW9/gNNqD5J+KKZ+/loqJei
mq3987cTHhNk7pORoGOy2sgM/s/kxJ8rLLPQtULrf+iuhiiuM2XCboHrFn/cKAGAeocjOgEIBgSV
of2OhTC7zgMtNXAMphB1qAAbNk9Lj8jXs11SlrvDRfIotNKz0JKjRMjT+Mcn8KDzVzQHdAL6ZoVr
CH/VDxBK29b9XeC4n7WHqy+k+4QrSR0K46Hj6/eEq91MD5vtj5Zm8JlZnGjjF8m26IGJWIOpUNml
mHMDd/0EB44YINRDCr+5wNa5vuEli6AaxlcCLMws0JNupJ/kzcjaDRk46EQMPjq7lTMXG7sptRJA
H2uWyY5OD2q0hfx5UKiwh3P8MuCDKYiTysbDEBIkU983VfGpseGl2iYQ7hMpuXa3+rr48pys74+T
HMbOWTWTekQ1eegdRS06RU2eSDkzLhCKCo/Z4b+bVOblJFjxu0SMrsAyQJgeDnNMT21bc4+TTvbf
leVh866v2RSVy8XoprdXp471lgWUV0pu0gX6lf5kvnjTGA9ubBGdUYdTHUCyKFAPCijnO3g/TRB0
6fpI3o5eLZniMzwwss1anX6vWGhZoNFCjZtZLjX3dk4r8rAAqTnKYC0p9idXRcqde2QdfhdQzcdu
mNc0BuUf7iqx69nXwWHB0RwviRdQdt3EwyhsVwbWQpU43GChWaY/0KprIrOrM4x8Nqr/sqxt80Po
Y6bN73C/ap4nHpwOWBFehCDnxWF0vW3oYn9YWSkDMNebvwFQWVXUiymkei3cRLCkiKtp2YsrzyTJ
6e2SFMgVnLKRfB+os9PkSz5xbRV8w1m3VAzdxLFbnGLh6/Dd+R8LmivnSPRZjvhbbY0huSutUIff
W2P3jBOedt7y1qMvRGlmA5I6tS5GOzurgjHl3cTOOh6nsjzQNVfNuOfq8g3pRQIwX+/C0FAJ/n0N
mJvBxqglXTsaAoeFw3zgEVX1/IYgMesPnHtZBJQfDE9R12LhxmAyCJW0ST+MX2p5z7Xx3P3WbFAT
+jO4t9PwksN8EbnevUPTbie7eVSdRn4a0bX7R9FD85IX1v1xuo9p1gpcNfc4ME28+Fg3moBgsyeI
0aBMdxFjdSzrxXr9y97yZN4G38sf7VubrJGEMvjT/eQdHIC1Yj5tI/udmxcNL2DXcZd08NE415N6
haKAKZU10WsNsTHb1Ndc9JF6+giQr70uH9aRtkRMQ1tYv6xmqW2Te10AAPIjP4o5o/rNFVLkRKmf
Ezt1MH5imhvnbu6o0Ue1YrWqzFTcX+kGTuRv1UIfT8kUGyTTpz6eZ3qxx48dyTIGdRUs6SuYJW6p
SQ5fhwyAedordAek46OQX6DGgQ5XxMMvqewY8wKjG1i9BuvJ6SBkeGYcnJgf4xBt02p2kwr+tTTC
40uotY03m8UaTRmgdrmVqsY1Tpb3zmt7NiVPdYzyp3B2R+piSJtuNFKnQQcMjqayqbd+lcDVefaJ
YL34CEKV4tkvoaSociA54uZOlrCprvkFIMf/f+Mc9DviFgEUO29F11ofscqUSJegZ3CtJb/XDJM8
3BdcCA29KzD5vWLaUB2ccLcuF0vo/RPkDEeiapekGgW6xDPBjhD6tT/ZDLE0sUOROtpr/dkH+6Q2
V5X8QrkaKF2+rTnrsCLP2QhLgyQOTS+6MC1dMZqkhQ/BzHZyqUFUjhzZHHspEQ3xbcPhsaXaPEor
3vScrTxzO4og7ehRlcnoRIFjct5blYGC79QNHxlkclXfWHDHUuTHhvqwZip+VCm1YS7dMuKy6e9W
Zz0RA0oPi5bp3GkYtEFKa8VOydJtCpOoRBTnzduvl6h8MtiUWRJVuHvm5kd7X2Y1aED6dIREKp9J
iM6ezh3gCFXljfW5KhExWXify6mcWemkfaQ+PFedx8ChC0mdxsFOHqmZLJhYPCD2Hu/nE1aU1B+S
V0QZ1Tax2NPl1+yQzA/70VsMYuutD2U56JtSl4Mowgv6wGMWahPuHhbRdeCllPIeaOvGWYA66xaO
Fjr1wbKg2+7xlcW9VVPC5jjSMAeTiXJTPSwRVqqIjQw20PoRoqPzHTrJ6qI/mKC4ZRWDflu7EVah
P+7eYmIDPCq7DRrBxChiQj5e/0A99q6FY72QH8SOK2A/MvJTGqrshXMTL3xRg/C1fcgyyBDaWTpp
zSyiric2out7/haDAjPBQ0TGahpHdomZrk9Uo33goiVLDU3K4bxYDpRN1KDFOxQWP9pZmFmuBygu
AQq49elc6wUuaA0FdpUv/y/+fDSf/p4F8ur3OyXO/ktayK0Xjd4svQWvep0r3zDFW+TBgc+Z8rQv
2xNob3L2Z8uUoKpWfDqFKnHDgkoMl2e8mkLy6FqHJ3G0S1d9BZXB4prC44/KdVy81qQqiH4rbc+V
FK02WHXXlc1cr3OI+zSkg1caLCwRywfZcq1wK4DtDRfWVkkyFSc7nCbQGo1W9Oo+1IzpE6T0fxi4
BtkhPh6oGycGcCEFw8/v5oAaRUjIT7FJ70FEUqjS59mau/cBgFb3RQg3uWyfGp6dwglfCJm1mz5L
lEGUEEyiAnqWsoE8od4+bewvK0VS/KYyPPuk0R04QAHOIO5qVsKfcKAEnmHKLeD1FL+n5bcuiVPu
JoYr+MLDr0iDTJ9ZWo67qsHjhniKrE1LEkRPf9hsO/48scJoPlLGJKBy/x4k1o0SMfc6ImImZkr0
tihhjPbVh+wuznPoFh3HTBiPT0VBze4TM/2X4IdgsymDb/1O5Suc8V5cEkhLYUrEBsh7h9S6ucTx
VAWqeOYsgRXJBHTNEyJ+qZSUlOsvKwDollBt/KE6n6zb0jM1tV/Lzvo8XnDCeoTJEUnSR+1Cpvf5
yjc+F/mElO+RxeKaKWzymhX6r9vPgR1E0ybBoxToopgxRUkOI4ZXi/etkCiDKC6cfs+PJKF/hKAc
ddrzmgW51ovuO11JwKIridUG8OPmqqR7uvaeEQZXI4Qbi++1QGZqHvCV05tBOCAMS6jkEOOXMwTO
mmo+QsAVkiiSxqbkjvSwONZEMhMMaCnUpufkTBplT2KfkdIejx8KZhJyYCnawxJg006bGf70fbb3
gqrRB8T1sF2hXqwb4OL/bEcroRmevNMOniZqyafmfUKaMIticp3eFwH6GfFv3Ey2cNF/kh5rr6s+
s+ksccSR9PXljqHdFh9vE7DM+lsuhO/pVjUMd3G2fjTNWGXJ162TV7nSDUSw10ad2QBz8B34gQ4h
VQe04Q6pb5GATSswdWrnmh/VpSnH6fVYKZr0nO7UivcLDJvVliGXDyHofBtxVt2D1AMWrsyo/b7S
j3LstLS4ArcuAiy8CYjbCjAmDuD6jzCcnx7fdq97MglekUBjqCzO/N+4e4U8MeDvBplYtQ2CsXL9
tVrhNuB1SaDO+zqKjSZNGw5lbE5XFbI2hxppsCBemLaWNK7s7KyqELOm6JqdUHTZBTs6pGZkXQ+8
T9PKeC9SdjqeIH/guhKzFxIpElWgwt1/RCxZ6WHz5YD3oJed2c3XtoE0pATEsg77BdblYqAiHNnE
WG7OBuWmfI84J+slEoN+MPWiHvVlWyuvyudUq7ozhsnM5Y8xsYNGU1532YbZR4bMH7Q1stmmAyXt
dijVD8NY2IFS+8cr9t4bVITxepfBqOR6voWi1D0U4mwMrBJT3tUAXfbVWB6M+GZuFeW57gKRQALt
0iknLXl3QVHB5JKMsho2T7rWL2bkZaBzeStz/F7d/Q38M22dm4G0H+rWRycZxgZsTlRdqBSt91TR
tlcOi0BKVAIEOo4eyU6/2Js5W0bDdQT9YPU/TN+Ks2nfyKxQB23B21PyfC6pzEW+uMVF5NZMxb1s
+3lVm2bblNUVI4Y0oO+Me69KJ+9vF7nGezgx0NiwiUsXaliAEduQY1qpZgVqgULiDer88Dw98qOA
+gIpf+pEY5mMwZZLUQ47JaHf16H6qVAJ0znLZDGvoUvaWtepWXMl137NRO1Eb6ZpHlwI145erj5X
V46NjLaX19HukuU4wltKf6c5J3NhrgxrcrXRo4OFHsEwbC04wFoTsvXa3kz7BVo9nvFGBp8Bxh8u
CfjHb8oq9vRon2Bi1IZfdLEgOK/Mo/JjMmzhxe8F9cCA6m9tZUFfb58naEz9zXbmmxp1KcGBX3mB
iPYc6juY4Ii8wNQ7cxf3M6h5ik16lbkiFasrKvhdjax5x2XAHt3eoB8X47P+LlvQjk4dSXEoODNj
w1lAcr5zlKoNq/BGLMvYNIBovP9nSDEk1548mT5Wzpkp4XqAAY2/OCTBWf38TQ0vUDZADZRWxCLw
STQ0OPdx6i1bHA+kJAqcUXmIJRPguFaFd71+0f62aRQYEaXjiBVS5ugTIVrlcug433HNJ4GrF2fK
vFKGkcw+SARiOX5F/npUwvVOQ6aTHmNdqyHPelzwrk+Yas/AbsWY2Y96AYixHCtXpBjfIywwWDQC
prSrc328NIsz4mW0U3+mQAKgKsS0HPe+iRGhM7zoatUVMJjvFOalT/WBp6j+5hEdOpMlNv1+Js+U
wf7BmlOPreifjWCS/CcPv3St2OZYHBV/RUmfYR8ieiCMPfqntSh2mqjFfgKTzCm0kFgIKZGafyK7
srEOeG/t3Yj0GFUuBXSKyOniUCXnlDBu4M2KKsRq4JsipsYqrLNFjH7i8rXpVb6Vsn2uP6ltA0zV
42kXVSsK+U0Vuy2pRPeY7z8iUVCcx6N+m9+wTvpqj8ouSMPL7B6lN88tyExQ0/RPuZcX95cLaMrD
vfhYR29RWA6/4KDCoJm82TdydgqfUlWXkWPF4o17irFfsqudYlFBUUWoYYSm5ExhIhMDpXytZa4x
ZhLhDKxhGk2Ah4kL5Ow8ESwGsJNR4LstVaDm9oRnRCYHIgizdzs15NL/l397HbrNfPSkk8thQYXQ
GKvFhc0gYcIvWUJiYrEO4YnhXPLqPJrJChouSCfGi7K8V10kzX3EUb8aWZd4ws8JD1WdCg2o+17+
C7tm+KSnhv6Ut6Y/FsFmeuokGR9aLs0K6whwV2O0QRzKTuYPUfPPoHAgqwlaOO7dcLhr/9YtGDNX
SmOhJu8xO5AkzaZaCayAOO0DXsWr0eefXjZnP7X10DOPH4kwQgaqa6tSfdjh9btpwClGrqj1ux5W
ouE36mTmP+LFJk5R3tsuhwobiJm1pFr5hKxo4eANrIFmkcxzhsKoAWvm/tCOGltVpIZwNkRvhdRc
mS9k3pKrYX1ap9p1NztnbpaFMOPlU2Yah50N5iDSRaraKA0nwSXI6wXSZHjgBTSGIV+7sum80ktt
eXC4XUci9ggxuXWBXdIUT6umjI9H9I6SYL+nAWKP2Sbma2W3sS1ZY0XneCFjGz4vpJz8evvILXKV
f41KlvF2Z9EfD5TQRuqiMkOgX86ozCM7mXeoTfhxJx4eepM6rr5143/oXfo+Ao0n488qkUJjJ+69
wob5pxOTMT4QuiiUZMp6bGeXP+l7BGpbPWTE6067Gp1MRnQNklODmqk6Nnk/7ATSk4+bglfN3cTb
rycGNvhLeM6ycmajCypAb6HtokXoxRKn8WbZGQvevmq6ZCHKi6hLbill7YuxrbIYDZbSpvBHH9/v
lKcmFndfJJ1Ev/MOlMSkW2bY8N7IkE5u9QFlHvoiwQbFYlMsgcln5asQeYTZ6LmpvYd4nw+KwlVE
xakVfs4HRDOhRJKi7usHoJRnghOmydRVGoHKKusjCyWZt1xi1hOQyzbUo75tygmOXmevBO59qw2z
XqIfjFIluqfaq/XIfMdVmu3/lxzlnHggRvaAHrHkDAH3nRIqjsNmvJKBUaoIhRiaMx/gofbRfCuX
NKt1ezsvJsyi2eEUCRjX33WP1cL8QSF+NCFvTXe7+hzuPPQIfMGNglHXTex1rR7NOVHmlnzDAzPr
+7tjhkmGdAlQE+KusQGl8bNZtVSN/2d+wRjuusTKN8RnRlgaFWiYRPEWkAJmTZhN9zY6byQojYS1
a2BqMaEztuShF8/lTcbgMCw1soyUb7goIVAlYCaTu6+pqt9V/EcKHYsvvlOPytzWakqCP3b/SimX
DwF9fSARZTvnFH3WPlF6btCEcD2DEWK/hA2hogfkvMHVBPOw1chAiecMJGPSHYKSZn0dfTJDgDMp
8c3fcKFFKchyHthMPoOp+cGS72FaRYqDJzsUcaF+XZ5qQd3jMWxZKsce3AyFhuLo34wMB38cpaOw
2X1yc4d3C9n1haIT1BX5jYR2/YoEWhVMcn2sXuaF0HwjMzj+klrJWyIoFM7KguUA+K/nE4aoSA6D
knwVSzXQmaSN54h+PJ/pymDEdv9CBNiQc7E1K6UoAZU6M4aAinooQCDgJaGT1RN8q5jUWc8b9dJW
7wIQbGPajAHx0UNKXBk7hHNEsLvW8J7XtPouzhx+tlUWqVvml0dWcvbdqdbK3//pLwQxjKp3FbKI
V4xWoZBbYzABa7fo+UsAnwI/bmQsNHJFm7WljbetZ52kbmqLWMjODgA0G2UQowrPcSaXtpfW2GfO
gZ2RZzMXSY9wWBYzQPFmebK8UcVt6A/MBJuuO5NH8IoflE0FEfP5na+UQHpYNi8L/ljJGwH/y/cw
STpS1uOfNnTGGA70RyVnvHa9nZbOTWVQ1WDppRt4Qk5uTN1EBb7L5hQ1d9OcZRNdwcZmjYEff/1Q
9AL6FVMSSD4IsXpHGQl7iD6foFic0oEx+YBpH1yzGNCyoZIinH5q6kFtexpph5rVc6LpBXpo1hYB
QH3gW47rJLY9ecsU4yWfyT5dnFtgaKVWZ+29817hEdm4dG7+VJkoRhbtFKhX87ZmCZKWDShAYr6y
ag5FC0LLEKKcTTbGBwv2JmKUNV2ZS4wc7IKEufiXfjc7BQoNyRTVtUtiG5JO9Dto42cYbSSoHRZO
vLuQiPX2G/tdMW/hzLOU6OzdM0ozJA2rQyviBEGFtaB09DFsC9tq+AVEtl/rw+y5HnmDda2Xis+G
3vwpHAluseXAeZdPYBM+0K6FQcWoTdWJYWi+ii2uxgHqp1azTS/q+WuPwVq58giEAAHhNseWQfnZ
IPW+aOU3ARPMhZij2+WIssehgZRKbGwVLpjxnoVzefeCurmLKqs7nVkMh/UuuAkBmvPm19VjqMkD
J9CjTCtYQlZHUze4DG4WbKWgGiZjsxNi7s3cWwvhTeEIq5TVb/9gUxBZF39gxoJwVwY1YeOrDP3w
X1dGm6N+1fHPwa4tYUwzKK6tNqqxSZE4hlvNTop2kXecNAqd9g5AvvGGY510edAIQRE16y6qewES
9OYiEaaxD2ZnziCnNYipFv+wZ/MJo4nr52y0oMyi15c0huY4w9SdUcPsjfioJjCe9jXC+laVesrv
n2D342Jj0rJHOas69aG4vci8nVdzJWrSvkpY/+me7nBWU1GvJA/w4+MHyPmCbc/g6r02NjfncQo1
7o5Rl7rmIWTDJo2w3aphgxBSMiqZHZe/SAGOMaQ73ovWp5LOCjSBCur7+PkmmNmXiz+nFfFCGGWn
4zp8pqLbiseTWXXXTB6cSnEUkG2OpoXKLwzdXQMFH6TOQjj72D0zSwIdhrhwc8ceRBTL6Ko1jjt2
JJs3gZx9Ya/hPzY/ylZkZ2exTZdV754WeQFr5/X7AzAxkzE2T4tzDmLxOe4AYQeOcBdUUZwqMdUu
8J0xvJ3ryuXT7TcU9w4/S+JhftY/YOVIayNANRNwMCfNBVf4SBAAkIm4POV/Kp7Ut2T+zcoKC+ZQ
5T2v6Qcy1ufl/kkcOCKS8yBcpLV70hIjMn/jfi0Iy0QhMyprbpXg22yIxYArjg1U7WfJvQzkW0uw
LpPdnYIKaSP8q43owiJk8hsQc6Pt8Pv1WcxSb5VwqgKZ08lqEFD4NNhDSRcSyIJFAy3Du4UO/4im
AdxcbhHt17nDYCyvbA6/UCJ/IbYcMAnpAtLWgBC/LaH6juXM0Xw/6uP+B9IBW9XDl5ybF+DBNtYL
mbMDlp4MjnIk5xLBAqDeXQ9l3nhSdvclh2JinNxUZdi7VdAexUF8z8qXg0I/a9hG1JIBC7M6hjn0
0WwmgFooEmiNex/S3Ntxu7L5+mqIDScOofiAHx7znpQf/6wGhQaIW3qtiemNcyxJaCZbH/b472Eb
s0Z8jLQFmgOxhWBpHcuDpSLZwzixbjw8tB9RAyAP6M8MVmZtff3IOqZHmQQt8PvJFP3JKYyqAOL/
YpGmS2r4oQBykBREfXyIiWFx1TQRZlIge0AbTyBlByWs2cbKnWDpbirvbm2gsRx8gHrh7KRx5Ibf
NBooAl4P5NDYH+4GqYcUd4USK9lMqREplSFiUUaZoWqgcPfZ+NZtaxyzJbE7YDJm92vJPjvwa3G5
VhHzxcGni3vniZwR2IsNZO6u4ySJKVgjUvzdGIILUAdCQpB2AWtDlQtrNda04A33/x0JHpNo1GLL
WtVGKZmcm3EIKAhDV0cxCqNR0ac+Rnsh0h3+hfHrO+P16hrLDpGD08mVsANiZM0aPLWww0AgtAep
8CDXSh6LcORz3FU72ur85GYd9+mlGz2RTLgr8cvAF/Ps3fKFTzLuqhbfxVgi0aK6kBIbnUYaK/BS
g+Tmsa5uqksDsw57a1k8sgSZ/Opp95TQCKgeQPqNXvInonN7kGA/uXv+pPsAKnhP5668ozZcvwCM
Pne3obHJAYY/LeZLrO/1HKUXqx1+XYH+ekf+GBZPrAl5x6PtgzfWfB7wr4ubcE4sI/4c4El+z5BX
p3x1vh/GKS7yK4+wHF9jW+G+uF1M5BHrB3PKDgUEf1ocwbLJor5GvSp1OFL+GUanmvN1uDuSQxtT
SL9DeNxoI5y9sz6up+R/X/JJ4nIjkKyqkOXzUsOrFkCSM+Myr9pF8+qiCiCddwu4iybLM3F4d6jD
D0L1zljXjUJ6/KPnp+Ry8muy2yRWfP4zXRLQUgvOStqNlFoW9fjKf7082eUysn0I2oJUXQ8Yzos/
cdhHoiGUcPzxlJGV6vsC/YiCjVcmDzTlwDi5x5TlMpI+o3XIlhej+04mafMdR8ReiUnznIXFvyth
V+b7S+MkIgRKqlZh/0YDwaBpM262oDeHyO2CkuXXjlaBCLiSmANGLo6vbMQMOY1ldd2KDHKYVsvf
6mVUwLbdihk+w0WDuCw8Qa3COgxBmTtIrR6E1spLMvz1GZY3QKN7onsx6RaD7FkGUtCunEg70pPG
hMdQ6F51NKn+AuZJ+Uju0reNfjN2SmsSl/63rJP5Rrb4MHWp+2WUnnZOBh0p8S/EzDuyXaQXVybn
sOZUzbW/hnBJ62dyv10SF6D+kd9fctfOv5GcVAxEpTd2Uvbm+cLDGupEzE+Ylxzv6c6ALuNvW6ha
hszjhBd27KzBK1y4v38o2eM7MhUkEZClaRyo6f34S/2ppR6sVKdHGdOrlC4xCO5tdFv0STidW0Cz
m+CuinJ3pflTmeqBL/5DzVbDjbXuJHKSThuiQUBnWHRwgmNlr7KZhrb14+QexDZdn9iPk680m8kX
2hf0/+AKFvs/ct7hCk5FigZn4c3s8TbG5+ulqwEBI2AbAFNOoDIzWBJl/lUWNn/feNjuxW2I1fQ3
kTt5iohv2ISDSbSvNCeVPefHePGOF9G0lRWF05aSNm87J3IDCL58e6TLz4rnASGQWzQefrCDCqZa
G4W0Djp1ZctfZR+Q3E4bnNMJf1aUHZAw8nj3NGu3fnz7PloBU0f/r3f0FawlEMHYOCf7xBXAWDdq
1ezsxAu1Dle3DQju2Sn2WoVcIpNNoqo1U9J3HEsbOKzNW7GLjaAgxx6H6y6zeaNCvWWUaLTTp81w
MTAUDDQltbbiP9UJsn875Q068uDaUj7Un0ZCXruGJoi8l0H+ApOyw8bkZ4TyBlUPr6oOO43o7Y5b
HEZ9xlVJJjd9w52F93zM/KwwvV+/xowUWu6PzzxSkCvdaW0TpgJWDxhVIS6eDsJpRAeqBn2hhMWz
tl5z+frLRtCybC+Bg6ZXtesmThAV8j+CkNl/3gBXTgmX+oTmvA8TnG5wltvcW/iLn34Xe4NyNMfj
V6g0FT7kLbrJGdiETKawdjlOgPxrUzMBmz6iUGVDeZyuKXTyYnhpC4SGob023KqT0HOEaSOHZ4KW
bw0KWWzxWwxZqTe7WuoCfNHexS1H63zfjDz/Vie+PX7K6WNPq1dt1XBMmfQxZGu57USldNNpHVAg
bbVVxpcYKZhN6B0SQyb4Cm/pwkvKe5tOIVjsLKom7yX47cbPt2Du4cGqv/cPSdLoYdiMmFuaPvP7
Lg530Fxha+6W4ED0SBuPvryGZIhKRPBF7pyfM/cqc29cnQnf7Y41K5D13lc2W4MCl2VIslazh+l+
pIy6cuMSou0FWIEnrSkW5xpCf7wb7A5tnfdQiQp1Z1tVK8FzeXs6LY04ZukNEQYtSm/eHaO6HsbN
Jc8Ea3GeRsNVB10g8vRqZU0hghswG+yxX5QzugESdjPCrFM173IjMjh8gBaRGT8EewisGv7UX1y7
FAfP8BHeQwVBnyHV42j7msC59bJbp9X/r5uSY3G2CVWNc9jXyQ7TPoT5Ip89LhM6PICuYFURycFL
8MgEoCeu9zt272dZm0rVi5ZA8MaJhUsx7S9JkgcTgT0Lw2M71vb8mGHhedPjPa/XHq3rLVCif6A2
G/i1gPw+bGNDZDvRtWQL7VbSkT1JI+AxGi1RuBm90dewF4jJi0sai37/+PWI/yan0PNIfHASjLdw
2DK01ajfiCqDh/fJ8aPD0wt+ZslljZYC7b82gZZ7cdGZacTe7bqy6MOgKlHl6S+XJN5QcCMvP+Pe
/5UOxREx1WucBACkVJwS4XU9eiF6WuJAAX0/Vz/dhs8iKYzSGXj/6JontSrTh5BG5kggYXEhPLAy
KGbuqVdcFxWQ8H8YRWCE6cI2cQ5W25X4zRBYY+WlOr2BPTrWv356aTK9TiR4IZojNABqC1p3ddeJ
ZD8emwR+K4v+g0SHXDEqtQyMP4dJ92/u5eWqiP3M9rCzx1l3FdLYqYQwwqwV5DiYKV6xs82KwkjC
GsE7SHe+ADsJkcYe7o62OfQM41b1OdSOUDDxq9MyxqAzGGX+kecvwm4o20X1CvSA5mqgDCL+ecv0
J8BUVKvwfUpy6e4zjjFbOyazHOqQp1JLbzQlpCGN7JYmFGnVr20xz3ogEPHiD0tWC4kDkpq/Isx1
P5wEzhHUthqC3o0koSPkQJItXp699T63oL69kFYJJq+8+QpAeb4c8zt77L4BuQdKbG6LXzXNPX6w
kzLaiKeq2/4qfwkuNF9OCU+q15Xs2aM4NjwDFMHxp/UfC5UuL6XN5k3OH/0/aa+hH3M2mif81+KV
sv3OmuGBwPxCh1jtARKbIuMtqt3lWhOcrP38vrAg3+RYbb9r5C1vA+DsmlvUJATsOSz7M7zLEH7m
CiOyxxYUSx2DgC8E0oloQj07R6EIcr3yqx7nIj/NVuv8xqJdLNN+HTN4zWk6arxCGvsA5oepxr7Y
e4bbM9xR2HshjCu+OSzgymqmvT7BEk3b/E2Qacm5pgrYM+LxiJnThQJJ0T+76+TJgMK7m94jBK6v
JEt7C6sCfEaqTAh/aqHV3HkGJ1+Km5Jvo32Z5Q3pb/2iF8RW2EqDvHb+l4Ol+qJWF17fXKXRrHrJ
Mj+tY830LbP/Q/hsje2PvdD4mH3c+0cA1eLGXBNrzA2kx8gkddWXHlj7InJdROdT4E4Sy3Sl417K
rJ0qvLaWu5FDiZtG39nF9bQBOT3L0XD3O/szDXb8TNPGK2jJgR2teW+vq90Izx78r81zAK9UQgxc
er2rRBbbFVKTuO6SiXqd46gsj9Zzkibjr7EAoy3O1C9addR/Tm/85vnoibY9ZzzotghfJ0nADbHr
Ml2P9iokwdeWnKHsMIZV0LxoqXcA09X4oaGfeexsblfgh+pGiJRPWycb+faZYnPxtoD4f0RsT0lk
Mzj3OOXN2aRZ5AbXluP8Dkf4Yf+ufELRyLOoIOZFSs6PJ4IPVcd8UCirL6rN5Zu/yjifbY8Hpi2m
4jBEpYhT0bZWj4tNGscazAzpOQQnJ45aOoe3uWnoxC6Ag5NlUy6V7WKQB2DbYGk8bbaqWWs05tdv
jATiEZe7BcbfdSKKXIeRmYk8muPsOylgZKybOvt6BplSvVNP13xsG9o2bXlDta9Y/WVkJ820+2kg
0HJx53qOR6iSnzBMZbuYakszjzo2Lue0YDDn3zj/cN1+J7NVYK7fiQnbOp/GZKxD8IniIk4qrxRZ
VpXXXg5jIQmQSjxmNFMOPeUxf3jq8wo0EOZMehci7Hbkj92udgYkrSqe3ZX88rEcpB9JU26TkC5N
6pQvQCvjlDgW1oT0LqnKwRSZrTQf1g6qWj7ajeFV6C9/Y3vS8C5UfnNvDVj2x32jB+EfTrfwNvAq
SQ0uASeHeJZgQmflNTjtRwWoUPvi2aA6a5xVp2DIJDc0ZPGhgFEawNPQNLPQUIR5GggBDitEo//T
EAg8IRuQ/J5QlpCSHR/f4rGLgqgztMKoGtkxW7jWYCfEqPBuwv+dLiWjyRpQQWtJg28sR7WuGCKW
Kp5G/tjKZ1Vkbjxvpu6j1fTcFVTezkEY33YhEy+ss0S8lNfBeM4rpLCGI5a6uUUn4lScwhMX0COT
UY9lkQb9taZxdR3BX+cHYro/qcSb19oExYlJAs9ppMDH5eGKvJP+GT1hfx8sP7SrmzLjd7dw0MZG
ISkZ+rPsjpE2YrOu9Fln+DEdqvM6TtVnLRsijzgS0fAkAa7mIS/GK0NkDisrK2a6d3RjIw5BMLJi
BdowBb9+yUAbZEnQ8ekfsYh2JrQA8mxmPessu/TUhU0HgLW3A0dhrSrG6VSMjEZURgZISl86XUTM
0OqHGuNfGduUQFAb9kJVE5KcAabX4DJP8d0QMe0TccsS/mn6NDRjcbZ8tqOIyYN7/cRySPhtiaJV
YHYkHyOs6kyXiy9DgoLjv/lFxQzVjdW1WVKG0am4QCZiQugUQ0SqGrlc4Xb7uyAKLa/fsAxmHWVF
xWDDLC9bbLiSWjSUWR7BeT9cJokAIyjhkbwZiivLLFXyeVQOtqWwuZrFTRRnFdcKGR9PIgM24aKN
q09hk4+oWtxQZmlbzVHwEe96ndZWmSJ91Lq9JDi65DWkAw4gN0M8AhDWIGt7UKgnjlFo1Ouzg7qc
6EMlJ29Zs2Mlp9eoYjxyz9K9u3d3HCGtjuqPlrirRwzeXDEIkStKb+YGSSDLrzA5Fpfr7h2dbr4u
auiqbWQvFAXjyc/F0e4LP2OIa1zm+3HCW8wBcTZ1J5vU4fcGcF1EK+a/blOlOwjkeAWPV6Q4bNOP
ipw/vFZ5uW8YiDlLsJMKrDOmq1iQsmEAAi3ZwqfYGhLH3MPVVXLHwP4vPgBYMAouucg7omySSdzt
aDn5OCXVJxo7GIEoMWjq4pfP6BaWgTQONxyUmAxig45RKtXktwIfcfPL76LCsVrqosEAUoOrzt/f
703Venf8b/JQCUn2uVuvAKFKRKRq3WTz/nmAPLM+M68WSouFooAxn1RjJ8uZSJ/oIIJHDFxsDxvi
xTMQi8YmsTF7KjmLuoE1EieOZs914ZVeWa0NjNCvFTAT/5Oa8O58x2YyanO4LrEW+zYz7J4twkcm
vg46Has66QKpa/MPFJ9sxNSAKuk51KDf2YiXqu+GoS6ghfEqiVvmP/FHaseNN0ArKueZQCLH0PTz
VX4HQGd8kRIxI1UW3uq6zElVKb+i/9X/XD7gj6QmgZcfr8oT+Gn318hUpG3fFoqizhiTYQoB3FbN
w45wFPr/SJaOcrt/bZ9X9nYw7eTLEflB4+39kh7Wu+fNchHayxFR16dPrrIuU5ECR8NCrEQybFpA
UNg6trBIVlYQdFd7n3hflHnKZHaheZVjTE6QG9XRSPyI0It2wQQ1HVr11nKfD9AKLK0SAexqB7PN
Fze3msNVFrS/Nj4BMWiSlpj/Sx09j7wGSNg6YM81WgZYplaKEem3HGR9JPylpeItLBn4x+mWu/V3
WIDRIsiZwyyWgDubBuKLcjFqF8AJYOO2IPlIOiuenUbnFSeJIHloA5YqMZ6ah9FiQEKdbuQT0W+J
YTPdItQejHNrqJGnxRR67xC2qUQHqYOacOF72i8aWOfs9s2ScT1LEofzQhaMTL5ouGsez9S78Sup
wIwrT2Ydrz0lTYCdi5J2jhHzJAoXE7gDRSN+bIBZafJKNq3g+FSWpOLqAm5ems1kDs25Uz2TbyxD
exmI4FkbeQnkVpwrJbbb1mfstGfxVoMvc15kcvW36SLs69PMXAEQz9iwYYQmMeAo/9ez4AV3wgMA
nIWprnpV5/czjPe4sPN/0Dvdski7cBBvbGHnLTayJDo8w3VtGjPMcL1rBZaYrpG+B4CtWfc7eehp
BOuv22FmjaoN6o4JXlbBgTunSeUJfpEFCRiOp02bC6UI/twSFa/kQeNvqStRTACzmNtQBUUQGgKH
cCDUUsQ067SumgT2G3y8KFru3jGsFFMvutIEgN2Hsoc1baglT6rGj+fI8fcXq7PL1gtP7YDFsJDh
A/LUaULNDc5u1rtzEMujDDJxo/IfnqEKNQ+1oL/GdnFafcUN2ZuhSEsryk8wEEklbd/hWyLFJg5k
r9nM9bCc7BLNU70RRzTS1PhGUIIoiTEv4nrf7TfTvkHws4np31h8fQXrP4aFbuStM0I/GKsMwwam
2oG49ug90rz1sNC6GWvJjarDLEZErB4uEDr11caoC7DZ20AtbUH7Fov4Oxg5icH+uHG2zOMzO/qd
1GCa6+WBbjmqxQDxdvzYKZ5V/ye1Bm08D3TpBJKaVU8WRqldL5CCWeuit+i4Iz1UwG9qpJUTwDf7
KxLctV8YgMrSXyjOcfXu8g8p5XLkLFp+VKamAHxDkjLIUbkp8Ip0CHeNKk+FRSPRK9iE7NvKWk3N
WiEHGAw1WqFp34LbXyjyG6lL8IrbsFT8LZMy5Fleesmn6/gcToYoQsA/hIGMNT+t8UB0t5CdVZrp
WmqzlBZ6A7HaMOY2UBPuLsMCYXe1bhSf89IEoLGjId/UG6UdwGtHaJHg7DE7DB/ECMgo4ic1f/sk
KFHKFqQhnxMiKkAJ04UnO/jl5c7Mex4V1xou5ItdS+AJVpcqKaEGd3TwRrqOdNh04rJJwLxU01EG
pvZtZ/28IG4Twis2l/xKkepWPwz1q5PqnF2VnVj5XLNyB1wBI8tgdavC+3Uo1Q7HUjSdRprj5NqI
i8LFQKlT9vlBVrkoU9BhDeHjVKZZ0QqlyG9TTuPx2sXDexdzeVoGq0m8GSPi8L+dyX/NRcQpqRur
62cLo6GYScTi5oOhGadjRp+2kzalVybTRT/tUqRQhMkuGaRbitP3ItAySF4dupbIzGE3wpASrLuv
JcLlJNn2kFudYncbLeTmATSnKROceiPEA8yG/1FmCbO2Fjf5Zab2mCBqQy/Q/liN5hZ7FXFaxqzc
n3S+461kORyRrD6Xo7Q6D8NV3TfjlsgIOqVumtZ5JOC+nexFmg8pWKclZX2qjEFb5yki53WjwSbB
/IKX89yITqVZvwBUKh5lk6eJZ3C+7eeNqLuZaOTtfOU/QBj4eAUYuOCWmvrXb32soMM4AQUxkK88
FmNba9LrNZdBCwmuaYJ3Yjm8mLrCL75gYkom+mbv2ehGF+I6Qma/qRrsMYEK3lzrq/y3m7YAWdMH
oTpfyfxWqU1RQsfcQA/UN7sE2UJ9F+7pqO1UfJTCG824wl9GQI20eReiLWkzZwmbrGpkbWQiFOxx
FYjEi/+aHsKelaSqCs3ixx06iGzjFEJyfZFma3s4n0nMEa84fPYlCB7ngwBTzasV99M/K5KbsK6/
Qqp6WJCNbndGai/vtI5Vx5fDCdBsMsY7rJtwdLgrAV7PgHdgbBVbCohZNMwvcVI40gdvUPvL1M2h
kRx91Hco9iZ1f1BDaEYw82yogDm8/aGNp4DzQ7fi1AUtAXXuC9uigiR7/y1KOnkLRmQwQUrIczOe
xs1EmrNEboJ8ARueajAduoc8bLCXrN7l+FPKesG10Xk5f+ngTGHWYDTzOGAEs8RdI+aBZDOph4wA
BOQu3whtvDHt+W8LMSe2alNiYM+HR8OnMsYylwTXmXtfdTdxVnDJwPKOdWckA5o4EXpand6hPXZ4
99Y5Wl4DHD7PjmZjbDIQ4acBYaF0ZCCD74fKCpPlXrZevuuYhFVmyrJjIh3twaD20HuG3TRHRtNi
/d0t3/KVhH/WcI8fokCd/gxoFMZxQW3KmfOvoXX/djoxLAM+rpnWAFPJNp86NJVD3SObXYE02u8u
xvB2l+/tKncAgPq6RXoX/5I5tMJdCAPQJFdS6Nq2TRXLXUgYHQMkijkujSEFI4gTwz6I230B5o13
dGA0gEkWwYwdXOq+GiDzx6CRWp8iuBTEhMWGArRckDZoea/9g6go7Y4WMtcBMuejgBBfJlP3v7Eu
UF7iSBlgbSfQH66NiWhJP00wwv7FQQ21nXSulNJlIFKRcbUS5sOS9fBhbFILaEThKZNBA5kIk8DT
yFLNEUkFrXs/xLx3GPQD5QVwRDWq6KrT8KCEMO7TZ994kRCnBrEvhFXx9Q/G+7zlWFZK6w8tr6uf
YOsIOmp7KdufL9gZsjOVIxNDNOI+0iEvV/ZpXCpOOX3pJ5yb2lsb33xJAIi096+WlApqLml6T2yi
lhP1f9G6ydY+E/bbo1dqDiD/t1F9ieqBO32gBatQviIJNp2PqutEnjqjnPUhNrUw4S0PXqh04ChV
asKOmL4FAkKYkWAd+sy7BIq/i+ojbVQQrTg36TU66C3PXvKcKCApV39osnFN+QRgRsCY00YwFcao
EIgT90Ce//CQ0Sp7QwPyc6+xYC+tT0YDe+7thZUAj9ijmwZ1ZerZ6smvXSPIQzcammbrLSo4fxIg
flKpIFyHGzKq5LaNUmO/hO7RlmS4dTfUVbGxO+hELOw2yiZJd7dZzTLqwK9IMCxUtze03jl7OlDH
3TMvtHyHwIgcsQwnRh/sAeooJM6X2yWICdOYAIfWSQT4qP0vse3mGQKGmwu25JVpJIphBhk18/xK
SkjhevfuRuTLEvzEv3dKBm3lYI5NfrtB61cZpJmsfy8S4tJRb3cnUwY/sEUD4B6UO2/bAy7ARanq
RQ17k3rbe3ZM/V+shqaNfCD+a9KEsZ3g+kVgWst6ICZPI8Bi6PMbvTOzLBcbt8rAfJdp2Cle4qvb
DrniAlB2mY+piEXPfKYZ29Vr1h5YHLS1AIVEDX5gJOaCZHViTLXm1KoJq1h5bQL2WOIyHjZaL5Pu
MxW9+tlJmPteKfH0n/Nx32XGs61ifXQ8nnQ4LJe5Ltb9C8nc8ZmGatB+NvReOZLpYgivBhAreIEu
rhcd3gU/A4b2xZGK+CNl2SfpTRQODVo4KgmnuwB0UgT16uhfLlSJLLAZi3j2YYLQ3XbEMd3DD6lv
EVPwP5RHEVwUTvjVzKgucqiLYrRF5LBQMu1+qPt/iljqpi1aZ4M1mL2US5DVl4KeIdFqzMUMyJ+x
S1dsU7QzEp6Fgruc93tAZvvmWJ+LbB9NrKyaXav0s5OD6NmfvHzIQU8RI4K7sSCP2Cp4tdBwHflV
/M0JHkUCLvJyZgnadMzTnXwO6EaoiHIYZILp0cTTAArNnfXBCkH7ueVxNo5L8g5DfpS0h65Hshyc
PZaNjpm0Afu09dTkQesv6eN34vlzOxaFiPQ9octVkg/D71jCv4DkduwItZkuuYpl5djeeJkQvzQM
k09+SY9qTMnLaO0TsjkbM89iGKoIdzApXzlvl9VfFUjBuxJahLqc49H8Rfq1cs6S3RjqUkLbx26M
Qx5NHskc9PqiWe0zBWEk/tlHzDSYGmNeGzboXzNl7YH0GOl76SbTrk+zFCibrFBImvTxVzNAktkG
DjNo26tQ7d6OQfgh2Wl2vSJ6orMbSDYD7oUVzEOUvazkOy4mgyy2C3kG09115AW2LdifAlyCGoOF
fX3NINH6P47xS8NghgbpF/esaZ13eSmdofPVuarj1RQc2GTxY01zKPdukOwhSf+KzWNT5xcR68LU
dQ5CikpJK8LRdk1E6qv1OdXjtf7G/KWgmpPFL9E9unebs/474ebX0mF7cYS6DR+HOVI1SgrOpErx
jnWurIJWzjVcSka2b6LVrmou5Zn2eHlRP0TiYqrkTWH8Ywn48NLWShJ/sxKG4tnjDA7l6xVxKlS1
fOhNsIqPrxofWh+hDlHGRhCJXPqoUzuKPD1YK/3LYpwpNqYKSVyo4G+VoILCYb2bQ7EUo6Q7F5PL
LKOwH6lQE0oA+QySHr5928Etek08FUX6dsDlASTKos2c8YN0KRohFbU2QDFeuw5RvZuMQuPAUOWz
UL4zFRZmmzB0b44Mv2SgDpp8FTCgo5/DdDaURY4FAIOXTZSxWbHraHA2nyuwzfR9C4LthG0VY4Kj
/ZspGSP5awm9W8HFtNEoOwEsGwagqNfG+9psCnWk30IgbUIofzbw6LLif5Gi20U3AtUooj9WBtSo
ftrhxBDwgM6AKqTTGQK2FdB1b+gTYOZ5SRQA942EI9QhiV+9T+13E5j3Gn35PXT7L47UauzjdFHq
FSa0fMmwD1SxxZ0emkMYVZxkV+HV6CRZ8sIkD4jGX9lAHUh6WfbTxM6VuzFdjwGNoJ452P4mOCqy
Zny1H4uVrV4MBxFqNNxX9E0AAqEC87igiA/6GL1pEoL/EU9H0T9C6nFuGB1lpDFRDtNSPIu+/Arg
daa9hR6OJ5NaNQ4+m4gGrbF4iGZ1zpo545/SHrCA9rokG3Sdxiw06NUwAsKYBu4VJFsxOq7ryhop
zuiHhfxufS+6F86vJThl4AYmqZwf43ZD4VdWLx/xJx4bWsXB8F9Wqh/h2qQLpUR9/r5VdW6e7Wpe
TN1o6eCRxxQXiSJVL1V/HjfnmUOVYCxjkXkiA0dIcMBMvGfCd+XDzbzPdzC20E+acrYieREX7SsF
lpfiv5tv+PQZJnSlBWxdlPmAK/hbiJG0zKKG8QIFMZIGSCfQA3UDJO1fTsELWNG9VWvYWCwFMBvV
tkzKu8rFgObfTOTg2nMe2V53jTzmIC9cfzjolCVWwYndDr9nXu4U5wei0MwAUsx3h/vseKXF4Ooo
2+/cRlSAhmXZeDiyrflFm8lnY3xyipiG1XByvJBOjz+wDhDVbsu+JT2qJqYGGhPGOVYGXItsLo8b
HbzRQZF0tPNNNriI6GRsZPD04n1zK4tgAdjCdwOA44xSc7jm0VqcERBWDcS2HJTZTho/bGAf80Pa
y/LKiPEyiRpYGQombXRZkO54TUhVAelZSLdU5PMXmebDJm8yHnaksGoHMjGktzQ/IvrCyWXh6vQs
QZoSZj2WTr1PNGtqjOb24b77oAi14DBoNoY5aDWwLPC4m0drIPu0SUrUYZ2vBhPXpNU0Kf7Su6l8
mwZ/RET4Kq5a1Xln0HktVV9siIk2g8KMCtccpnxZ3GUqNsiHZdsyAkBn6FyhbAypFLnSMe3qj1+T
9F+NU3zX7zPKZqofprL0nsvzIvzPBvqAV2BUGR6+TaXCxwy5ufl5ysgWRGKeJ8KG3ywkmPagY35G
0IYVUmuymkdDRDyNYnbJS0Zo25myAYLQUElK7FcqTC1yqCUGuO5WE3yD1uIv76L2y4WnaWt43dnN
5FyzmMc6pSqnXlzvSclh3JndOQHITh6h+Yqq7eDiSFEVx9s3/Fp0XzyToMr/mAPbG57VK3qkzdte
1roPELU/TVqtti65fO7ZynSXLk8HR2Y3oatuMazSDIsUwBB3kAc6abCiL910miM4tjkSEe4hLGz1
YbPZbsDsUnZvU10QOJd+WyJFKYbpgJuhqq2jUsgICAzY/qzsnI0PwJY0Z9Bnqfa7tnY4/6rtH50A
j/Q7reMmpUEa34EPjRjsynp7wqTXavdY/OEpQCfCQjKWWNR/S+4rDwedNiuXAR9VDNV8MFaGVbjB
KbA/78pjsRAAQgHqKIKFgHycse4ntFJXOjbwy/S9UFlTtjJzCL04JZ241nEV1Jlj9tid22P4lY2e
qhEpPTQcDrbgSd3t7v4WEaIoB8Uw89dI4yZZ+exadVKOP6eFw7fpFoYe2cX97liGA6jRjydlcUWH
RGP2QPjTGpvQWXMFU3nTsvw8SipijKy34AzxNhk9bsiBz+LDJ57ftOMWPbq8vSm3n9JYsZQFw+sf
pwhATBJ730/D6seNHmpHu1cxxc77ns7yg4lB+vPbKhR6ayB7yzbeV6wxlpdQcGCVEAEi3C46MT8u
TS1WSQ5G8YHmy5LUZvGBTblM93A6OU7AAy6DlNcGprloo0JUuCx4RxLe0+IzivNejmqpCBzU3eWA
eqkK5mZJCZV5oKooZw+YtvjbZ8rG8ZF0fhRDuN5cGSIQX56g5o1Mm5tAxcbGCxCSjcoX4e/7uhF5
fSh/DRfvVcy9moEbNUGI/UolF2CsEKqYN4hZfMz58XXKIqKXkxGR+L6eNkOBrTW6iDsQ+mE8Wlv2
uKEybOuZ5CAx4Zq05r5aM1HZASlHl7TA8p4RivYfKO9iC8XlAWUw+j8Mdn4DAHINPKxMu7nZRUBE
MeopFEdNBjc5JntQtJww+S4iCs5wz8jjjqu09ifAQMs69RedX1XdfVCY7D5HUgpq5qzLPPTBgfke
a1fgTpjaQxOOOFvOh6g/8LAMFOnvWY1HS8DKcjQPgZBCx+89oNJWIXZ35BUI2g8QymR/cDD8oOx1
5vXGPZhWjFuNalPBasVe95yOkyNJYD2rw8PeFAaY/s7e6zqA3mRoSjvH+8/mxDVdyyCyXQnf1R3v
nGjLSmME69yBHiNZmoLl03hh+NW0eeUYfxgiMHeU3x72O4qbQNfZ7NuaMyAecD1l4JdjiSYbc1iO
wT9wj6Wgz6Hosn071+NdjxyKzWt2vL71O2VhoxwvlnBoRDKpJLT6V283GEFNq8BMVKPd+yi45PoQ
Ibsr2mgmYZDB4wVaxGs18pZ/82i5O0bC2AWTgU8RNA64CQJewQ155XkBEx77qxUVGeRVxpV8uXqG
OwNFdU+UxvPCCA2Uwf3QYS2u1HGUzQk+q5Kb9zgHhgTjklCGVQdsnjS+wgtVu4QkUaZn4FRnyPR2
LutcMxJC92zNWVYlYHLZW1NLbhdWkNbgSrGJBuLgIZuDeBO0xIL+D9mKvtyIArxPJ1cXfS4G0xAH
rWiA62/BUUaLry1kMZEH3Q2YQaMcWgHH6joZrhknowJn72KcW7kdnc4UNMeKHBsHzib0cdgvdy7d
ymxivvSJ71Ixe9ho8nKNla+gJNTCLldypItjR65sJaJ37zwiRWh45NK9fyAev3BzT7tO1t1W6URr
I4ZGQrpDbcpnbGoCGgFPcOHG2yFDFmPqZhCJZUruCBfCepyeTMWwrn1MhQtEC6GvQXxkuGY07u/f
lMJ7tbeqbae+MeGY40mnqtHLHV7k6YtUgC2kUxqoBN2AcB/4+PpY4sfJJGTHlL1R90YfWfRZu0mO
0GEwbPLJLKq+M4LRsIY8c+k8W8r0OJOao4hwc1BLwTYyQXoEA6hW6TAP9naY8ciE0RCDGYuQVCDG
YuZJ/0YnT0qn5oaYy08onYUY8Ivru+mKrVkGUyVkOGXspbP23XsxGm1Xp77/ms6XdPoXV6Nzu1Ba
bOhBCMZgNXL1RPsgr3lWMQjVR5dgdsYw5AsH/PRMhBWo+iSgbY71smmpAExEzb1HTs93YSwni7OG
lb/+XJJwiR+byXrYe6e8XEo74a918bNfhjXwY8J8/dJyVKXfuXEDhdjgIXMl4zhoRibUz3p3MTjk
0X8hq7JL57wOcvpKyzB5MWjWcHaN7zbd22VoV/fHOycDUEIjAEZk7q1yFz/nNv8zpo8XTo2HcqGI
zIL4qi+d1feBDdihF9snQwRj+Fob5/+ZhQj67P/eyrobYFdz8FlGK1CpDxcXr7G6T4rlTyqiGx8l
sAR7xXUEaAgI5KF6gyaf98IpJmGY+OvjS7WUqAjylQjylSLfdj6N0T9swFemqLGQmTUqB98NmnqO
3uuoPR3KGQqqNe1HkedBYrjfc1n3vl+UI03obCsfszpH3TtVlFpy9gNXFiGZxVxO/Igg10nnZG5s
zSblofi6TiEmHJRtiw1qgXKFUKeWON277HFPfa1a6MoZ7rCub1uv443oQb2H4TUZz38nH1VGZ/Hh
XlDNu8u7mNaqxbhl09YBqyYZqQFhUa0cxeD8hu8bV/OLIp3Q2CSDmXf1MMxFjcg/jMrNcmWKyJPH
3H9ABU6U+lRm29bCO3UUgQhJ1F659tGxvq+B5t2CK5dAFJfQ4M03F8lE/N35+mBSVU0//7eoto8t
7YhJWg8SxCaXZE4T2jDFUEvTs5ICx30sqO59vmGyazWOD9l+AIfGGZm31JcjDyWRiStoWNXx+hGU
ssSqEOzR7+OGgvraKd6dM7da9RACJD/vzwTkESnDFncSWvfrjpXHNuZXL2iVzTMhxmp4dyHR7ZtQ
nUDylTdcx0jLiV5+/1m86QHrn0WneyR/oprzm0zNpB8bSh2g9wwpF4JtS31tyq6yHavw+bVR2bkD
SI2KRcPK30jdtj0a7TYyr3sTRU55pdLR8JQaf97Xv/yKRxZEHdXQmlgyTgWbQ/BjGeEBTcpNIytt
omHaCuUV7anewIaMOWav2TNZD3GbHbUb0hYSIJ1tvyqErhZ08wj9kIwtVx9ESNiKb8kxVxG3AUjJ
AS+uUrSpds8u/4rS1akx7XF6rD6OwTJEjjKlx4w0A3ZYj0g6hm6JpR/KvBCodic/RDwUuCnlwxY3
smuVmLX0wra9HNVSSsSTmtOr1gi5fCEHpK4BHN8oKmkJLnzuVdGTFrwNUVuvm93LcUkT6tyboq2f
2SYUT0HdJbTmdXHi+WNA4zuTcm1DqjOgTDbJ/8Cyub72LVz2KnXQeoUrqN29r5LVtnUH89wgRAcM
J/LmOr8udh1LplRyLW26Kob1gy5sGn74rZhqeCVki/g63c+x2MsRWHZydDZDzx9M1xs8bba0Cjrt
8hH4Bm9F8ZOKLebrz9olNBEwH9duK6/fSofEHtTRCBOYRGXv0jVZykUM+LaF8aqLlG86W8YzKnjz
/nLqBeFBK6qXuwFkd+yOPBgueM8usoi3W/LnNgIFT/A4LsnVi33PasHgyAFwxEWXTkbTP8U3qXTz
5djdHu3Xg4SmvN+OnAfceZrF1cIJlKqYWVces+VlJKAYOxAw16IyR3Q++FnLpB8lf/C+EPz2UAfv
BUv1OUBmydTKpMUt6Fq+mxlbrDMH5SErWVuuN1yw/ENexvFU9qZiEaQdrLCGguKlVYi1zwsjqEEN
mp9HhqE0ED8NSTM6ag9sDrU9A0mUnoOoJIY20THZsZoMKhN69F3hJb4ou9nLPPWScfpMAVBMQAbb
EK+QfJJMDNQl3jyq2F6InyyMY0cVRVPVMdHU5rQBkAZNfp7DblOWPK/nkLMVQ98yflFzMUK5Jnyl
OVkKUALLQjrAAjuwS/LEAla9PJn4s5S/eQSTckjPPLDzVl4PAgoed4s2y4flpyh71IvmMGtkP0C/
CtK8QWFF64smYfbms28EH1cKwAjPqP8+eQ2V9iQWvtoFHgBT62cjNp7Au0bcka3E0plTA29iCr1x
IVtUccyxr5/fPTU7vZ0f9GOqvoGo1Xstcn39Cq2zcKEhjsaZkvuUShiRByzZHWyMbe8FTbaJ0YVO
I6ZH8tPyqBh21puVMgGl9mdnv3IRO34PPhWJbaIyNpQ+B7wVs5ojg0+vVg5uoqg5fczsT95jk04D
aed4YHqViw6FqX1NUnMif7hJMktaJ97i/rx2FScQ/JCqKI0vPNKMCwkoR2IxTXiaNJDe9jNjC4E1
iFRcecCcsqHC4RSE00AfO3PS4UzUBJO3+QqZDNKVeimWDG3ti3sM0lxXEhYvG1BCdvk13fNKv7Js
FElOwILDHx5VTqZIHpy4Jdz81NBJX9tzmMASmI2mIepmRhJ3tqiaiSRlPNoNrqdeKf7DI4ynRf2J
68iqYPy7UgKW7l8YOGE5UM0E6W5BSucZVqIMNMAA3RXx/mLnNdYV9sSvabBccYioDwwQf2nsZHBt
8ej+3EOyTAouz4hir81X40O+vp/SJ828oIJhexEpEai0WiAaczPwrNXgRYIfQUHHxZ7CxRZwJLBb
9KRvFqjl1YeKzVbSCQKpPP/6+L1jFpjS4fzBTCQHsY20MZfFffpeAbQx8iO5mZPxxV98bU/ogx5l
sZ6G5PdWPHRDVmvRMSE2VzgRqRLWCHHTlTJGVXBt+YexZSzuKLvwV7GroFdVrgas0NG4BAUkdZ1I
dBEP2x32v31tONUlD5JpA0St0AO5dPEoUSlJ9A+FcLqoIeFNYt/i8hwckXmffgpdu8Pgp7a3WYug
Siw5l7jhmF976NEMu3C/JcsC1MsKNcaZ6NPtN/beym60uX5rUjYHeE3i0V5K7lUxWy4fvUndp3xs
8m47jrcNWMmHfWKJ+5zitJcVuHbD7LkcVPUsaRrKWgbOZeMxkfqO3fYI5Y5tRgGQY+i8V4T+vuQi
Kevf6y1Altz72YuZPbDfulH/txaJrjcxnsQl8v0rRe67QkzKqyA7wZlXUw3xMKzO2NT/bV+PwlH5
D0N+Zr954m+QIFQ+fmaLQlAjI52hdblqCLWMI3YACOUxZ4zR/GeZ/xyWFLfAh1DDFCSfTlMg+W4u
vebP6v4tcyoednYNCGD9IzJ/l/6M4aPna921tgqc2vAzvuYjZBWdh+PV3B7oZ+cxkxdBHk2iShkP
lyrPAGyrdYA9+RwATZQC3yXJd1ixEeY9M2exd1omQ5j5eaRbloSps8O1Vp02sJBxhAKEW1bKEctn
FG6dGD/2uCzKqAEHJgMayh7CvTuV4t1xitudoG92J9F0qr74NZQXO4tTUZfQa7ycbD9tpiwMMYVV
TjE/6nbgAohacXQR0T/W0J/60uBWo4FUY0M0MQdrgMzhnRwFmNjzxDdD2WmPszyrZG12uLZxjh7j
ZH0j7yO1p3ys5NnOGSLqXepPC+TjJaVXIyPmZ1ogrj4RPyVz1muzAWc6Lv/38RDnfUs2ig0vTnkr
6ambFrxie4z4wfD/vTxD1NVdqobIr86PXc6mpllQ4tmOMHEhU1OZR69oe2YhM6GZGe+u9auPcDgy
ygvKD01diudynvoZ8oKSEL5gg0QRBu+RBNaw5fOLqkbjYJ72biY6+GaULWevNpT4mRyBt8HyBS9Y
hLY2pgEPOrSqGNL5FEH44EFWlvk9aQNmmUrf8kQu7e3k8GaCtRKWMVB1D6tBGXH8xkuZjQ4jdMAy
Kye6izhauKsjgU4LbjXfyVNhY4eaqN46b1m22h/vE5K4L9TwYzD3aIZWdvF2Pr9RTWOzonj/qINS
RPJ7eAw2sye9A9l0k7yfHGRrnU+udf1uARG0V7r1HTHS1tOd+tLrTyNmibWMEJnW6umFpvj39eQ0
nYNx/0kbN/UgpmAOh2cU7EbGmhHoRcXMxtnJIkjZSPt40g/UEuYSBT8ixBfkjnQC9SWvd50exaqh
M5GQTPgad/torlpKwm6HXrkq3acHePwQB/1nFMhV615CT4N9/TinEKQU8JyMC8JviVWrSimjHgCl
7l88XuEL9GklXtnkrgQA6IdW0nk26WTbU7OfAbuNHKXJmcuc79bLHGglbhJYJYd+PD8RATOZ9JmZ
I6OgZf6yYQFf9z3FKDnKASxiRBSv2GxN4ukTw/CCl+uJ+Eh57ORFcR3uuFDseMO04LuYp1Vl/85B
MtxqJI2v9t4eucl5MHumH1Z3ICV9k+vb43HyjDKt9okJDZRhfzRBBf/hhNQ3qbwMqoE/Ixa8FZS8
kHgKlFWI9mSR2hjCCNCAi/xDp3spf0MzgiXVWXv+Vq6S5CWoe1a8vtEBtKYyhTZcpKywUU8oa0lw
azjyoC2aSHk6/V3TRKucTzTN9Jkw8uW1knjv2U1eJDtXgcbbJvfg4iryEU7mkQyLtUASuOwJtvd3
Hku4IP9ioeaYr4D/MAZE8HxQieGlGJZ+9Tg37udOr8IDwDBqGLrLOTeARMrTITrUinvcg9XGkhFb
UFHJ9e1tb9b/09bZUY96Na/H+yWmlpFKxQKWf3pdI9lUV0L0rjUxPtfpUn4fYWm5/hv9/OznzPMn
6JIqZ8LQzmb9RUhsnJA6Ma0BMf7lWUcGOZdUTjdARFePs7rebULEAlCbPn8G83zJEJyZbuz3NXyf
/EqFp/OkNG/O0yeyR1Li3dgTp4LvzZwLHQoz2+0xnM4a+BQZonpmhagV9RUsdpyDMDnv53dWR8vP
4uwW7gX++cZVd0MJlE4IdPPHNROIFiDxm5eTO3WQeS6ZZ2JX1bAX40AOsf37KNBymx16R30u/WX8
Aafey+FIrwaFmvyY6cyHoUbL0D73lWu3xnC0IIhRoR4b/jIwL4WtjFe14IPb97XKMx64jvNUSsBl
cGDXeISqER9YNbCMGe1ASA69gqBzDuz32/kagNkMO0uiOrd63Tq005z5Gbuh+ifDHXDmgT/FmSxi
tBh4tdo+pJCMJYfZaiwRuAuilZcixz4vTmfVIlgFEhz4l6JBH7GQoux2suthq6fol3sgOpUsr4zU
8IWcNzmUEazkZjR+Nz9fNgCSHpHWZjx+6+u7VyX/BOX/sCjyB0CGCi2EpoUApqac4xh6c7PMRcFY
qY7jyJOno5R5NuurhkcoleEUmrkTbVDYTK4W98WPWtNb4afG/Yob3T2cP3tDgHEs6e9SYQKcdE83
Wm09n4szWTKr59VAbMp3FUh/I4G04wmLyK+cS0edQKrZuQ9B/aMBoaFSOMtwrNsiPDZrxnyh8mYw
RTxH92jJk7Niphui7A5skavFOo0mFOak3nNFCu9Fu668xhENZFS6ifQT69L+seLPNW5iBlwfkO9l
OLXhfi0G4VS+oyaoyCV2RL75CYJHPyeIvz0yKwM9SQAl6AmAA4YOcu324IntSMlueF4Vg1usKVpP
9mnKt7bgqX4PYY0o3Ewu9JOIVBFmzlijEmBwyaqUW3cqFI55rvH3Moy9voDPMrm3tvhp03vqdWYJ
lKn8zYQ47zZTKbJcyNsPQhDePLlk3gcd9MAEFq3XF532tddf7MWKaGleJ7A2fzWaSECUDm6jwFpw
okifEHcjjClaS++bx1U0KT/xuPpo64EKbrz/uihLkGWUetjnh4Uim2zCOs4dusc5qpwXLM00pRMf
hcVIvR1tWr0R89pYwDXljoxsNfV68fvCIPUsAk1DC8eZHwr70N+5VqUuUv7MrneBWUCrvMzSxgPx
rQRIf8RgeUSTXas3TUcH6F09XeFgmgj5wlGUgyISkvCUYoWtfUXf12VQkE/ey3f7+ETSA8RK8LzM
jkST67ZYJnUCJ7rnjcwa+NQKIYfMaL0qDfUQJ+Y/Zus+i5hn9vGRJthA/J+/liKVJhLZxTaV6Idl
yWTGUoOcbFtxBby3rU2koLFbR9Rqvu2G93JkHpP5tVUedZj6mayfGWuR++UKu3yb8Gzj2PcPhKO8
I3lt2e3CaUvzdAeiXRMEDrc4fYwpvNmCxJqPMEiuGgkv0vayjYkHYVnMFBfWCsQPZOgyvJj4R0yp
yAbgrbJj1I9j/U5WeFzYI02j7HBv70o2hc9sLd6iJqDYtGmN5yy4K7/n8A3fJjgas8263z2wfKdb
eFTRTFGDEp1jt0WhXXYUeJj7rby88AQWpjaXxo9cKB3pVYgu8GFB/c3Mso9o10wMgmZXOQS9PSda
G/xfXbp3kQWj3UputAdVSGcbIGVpdYzH9xpOOgzk20+vK2ce5+Y0Zqq8OGhD4oluSSQJkkd1oe8k
gDTh5NLl9XIXst0dD3BpuZqsRyx4ZzitybLUUaJTObuANzWIX6VmE7ZxS5e4OCuGyudAl9pabfaa
9gKXmqtfGsIHh0gqbvWMcpRioaFaQa1EwAbBmBFiZ1Jn8DDz4N2IMx1CrR3AldMtfI9EJ879Af5u
/9fuVOeG9vHcuQeVODHWqFhgmqYI7wQBvC6stVD74KXgAda7Weo8NP38xdX4DqQiG032rl6wa7iI
A3mXnRrGpgRiVCaKoP82zDRqb6fMd5AC66Ig+DA4DW36IMLapsJE3iBZvppzeQ2yCbaacaZ1wb+B
amWSX1VB9BYTbf+SnNGf80Jgv76Tzpumck+zQ9gSsWffIdoCtWmhyy2eVADjyrSmyeep37QhBz4p
iPgFsfc/BhpmqLYdmbnJ6yaziwztSbgF415ECXrRXUD1sQgtcUBBoAkurgyZbPjhCQvEhoqpLjrB
ULtrFtvyNE+TM/dN1bD866ys68lVkXlPXB0il4HOOYdUPSxwnGRs/BcObMU6ASgteYCwG/OQBW75
YmoYVdFqgQIUwjvsxjbxcB+JXBf04stMNZ1j464EOmSOevxpxedxpaDudHyNzfjdSDXe7wwlZ7ZH
X/d1E90C6Vg65d/gZ9sz9R4eH7Zuv3v3Tj2wQZRPGzn++zv6WIBPJ2FbjaQHvPHlRX03yJeTd1aw
Co7Weu688MBYhT7nbPmZ1Oko+14QQsI8N0uKHQeV+r7pb21TYB1w6gdgn7MEs8KplQSORK8LjttO
fzixB6Q4nhr+hQ3sdeZRXsmXuLCyKCOrnlSkS/76y5OgMLfDTcKrh4X4/y7dOGdqCovoreQmGVo+
H/+FZA3a7WqTyXgE54lHNMyqVGkFff0VF8AagPVdM41kDIWCimNu+iMHkdL43htmpVo3AnYwO0c/
Z+ZNO8L1pSXmr5xJHEY78DSGN8esRTN5Y1pZ0xi/+W9lv4tyglQVaTvGuN4BkQGODt0lco8Svkww
vcRkWNwY28jk3tOyetG/vjK6PNAAf0zzSub+leKDqC4OcT1eW3W9ExegjOnR7qOiY5lfFv+0LaTb
dsqG+M6WjmLomgd6Wd0yzB01r5oRo8zpZOXIR8KzWau3PesmtPWadz0JdTSUbrDIY9VZ64XA2o4I
Qqo0PVm+oOpTKJAV7FuvHsyUH9v6zyVhofe2z+uVU593VZYul9aq8lUwH0CqmDUkiEzqKdJRPauR
CvUgAMXvOPAHmApvS8ZDwiR01rzjQ7H4Z+zUN2aIUZCU09E+dvTSHVZfinl1g0fqlOhb7ekv6ZMR
y0yMiuGBj3GNlIn6oxoq+lZe3xZ5D5PTd9wixnJm4IiygRQp2OtOzM6Ry/MspOP8hNfrjeAAV/GE
/Oog0opYrWfd5h77SCxHrpiGwOmGvSw0zng6RkRnWnttdykWliXYPxQfGPBZwK4r9dM6kIOpfZZ0
o+MUshp3Ytr4JwDTqNQuMr6FjCTIidvfySP+W/XV1iQvOUCxZL8W/AhJwtxyWJcqCXakC7v652aj
INdDJQqi8qtYOnEbgOlsEPJAKpoR5oO5WdFbMWQ17JzJVDukzS1AK+M9exNC9mxfdNTTymUSy9OI
StZL9Xq1PsuqZe90JkTcDG7YAB5TBsSi5PQftbgyd3ZIn0j9yTML/1hQZBDOYty2dl6zL5ebf39K
zFx79tj7BTYYTKTrWYGvVMGLDAeEEE+hqHsxawtCxYvwWR+SRIkmddt3u1wVeqHf1/LNFeAORpUc
c8GYetwnU988Dcrjjpfn1921r3NI1Svh753L2I7UAf9Mv1qzvTLj97Wqf40UHFSXbbO3hB6LoW4Q
RugjmJ0XWOFxhG9RDHXtGtWyYrRI9087BKKgEa3xkHxCyTm2rXb4Qqp+QMo3G8pUzGmN98MA0JQH
9qrP1/wF52YyRi4c/3KuHROCI/DbRBSxTRU4d1savxGJ8M+Y2h60EAJH3N0F3WyEl3h8LrzlL39o
hdkLAbFgN1+zQoyXD7xWgifU88bgbLPkSZZaRwqThyyqraopinmumlwS5aqfarP3enrYenPC8a3b
1Hk6Y5BQS6zOUyDli1VCKoUh0XqoWIFNJ+Tfjo5MGDfuTUfegpMCtqof2Q8z26SgWOj7Nbm5s0FC
Mh2PwJ6YBw1tB/bFcerTroKyWfrvI/FeR78yKTBo38wYFnEp/1bErzNdWN5aCyxz5P4PrpVmuT3d
nw1E1v/MHzezzcTgbM7OU2WtRgvguH5UoE1gAyumZCpyENgKOlO9VmDdctv0B1WHhh1VSYZOoE3b
E3ZirzzRPyl2EI5zh9oN2RsyD/eVIG+LWDaZkhcda0ueaAPCPz5ijPfJDQ1U4mYi4gSSEn7Y9MzB
0Y7An7iuVg47GBTQ9v+JUqa7Mwu7oWFRJPYc16QZnnnvLSQuCUNSXq80fO2B7CZYkpV4CO2PmIWI
dR/4vKOymNEKTEhP0wSTuAAyLj4isENpFKhjelRHiaW12nB0/GUrilkVXvJ7FbpD4eI7GXgBRALL
oGyTpMN6A5LlWftub7g12V5obO0QyLAPFmOwnx8PtEx0L4Him+ECQm/x8T5esNLodx3QMwfzkj47
nepckGN2Eyb3pjB12klE6MYeTqvqadgyUQAMWxK+HcLN9tMBhfCTi0MnjSVhw4K5dxML4A/pgDea
luCNZ6WCdyGpqo1OQNR6JdIjMYgbDgjA1rmaWPhAguAxXEljQZ6cqZykifBZyM3G1F5vTbvzn5AO
D0VozQRtdGgrXCIBJomZ7eJTACYji+aXUeHDzK/+7m8ptVooDjvj23qgBVTT2dSlRzeWQf4zAwsw
YbjRHUIJ2tKp1D3sZ/6Lw3txnqrSWpihtxPbjbm1C3nhTdudUZfI8/gRDWR4h9js/OMEYBz40lZu
Ozvs8NrAFU37vfDnOi+gwrNEuDs8HgfEN5y2d/ZYaA8isNcBKi8mOz8fVE4slm+Njymw2jFqFEzg
ZFvExGdxTfBBJXb5tnO/L+tH5o8+ucK0Fajchc9dQngAf6W8662/ObMYH19ptyrOoPrvzG3p3T0s
9lorMpfFJ1IVFF1fYhmZdecdF/6gm7WVP362n+YoWw+lL2akPGUcfxaFAuFdS8kOngbUsJ4tiPGi
q6qWl9eU92OdGbR4RT09OzMJv4wRs7jAR4ezstUvCCKgS7b6iodW3l8hyn0A5hSwTOU1yAwNcqr9
3kz7VHGE3U4iAar2yqY25QIKLNFeVFHpOQibHsnmHMSrG02Xi9f0yxEeOjj2pAwZqjLS7DCkyRJf
XrFRklIUmtRP26UrGeRpsZsTdKBeBBqp4UDEiaWVPywzvaO6K5lWHgDW0gwP/OQ6eYNMSfQCUdTE
s8UHvtPWT8UrcZepMH4BpZ0EkyNzaCCKnPA7HeGXxxbf79yyGKJb6a3gpsvCMe+9W50AEjsovM1c
1DenFahDeL8VpypSdrcMsnUYNTV2cQE0eQPmPwavD1HlT2MZX1dkX2/TO8sMbHTviyIQ1hbkWQuU
cyCWHh/ozJbWpuTAt30u3asRDCjI8pHya9Zj7lm3EisA6xz5tdxp2jfUHAffTfI3NTA/B2dhR0Cs
9gdArO9vgsAwFTwuS3CPGSZIedAUIZiPBLQnDQIBvKyZm3kU8rhBrXOtZoHuk7St4FsuWAgIKY6a
GhgjdjRIyJd+X8JzfEhI/wnhOX4TQW/biv/zJ+fJdEBmH13+iDR4INNidJ0t7qWuy06+NX0iCklC
kUwr3I7jkUTPwnpFPIs31nFD5kVKLeOQEydSEKfKxMK6Yk0rOW30oXrP8CIvxNZPgbPlKXV031DE
/9ovlNBHFpjCb6QdTw7FiJunKde6mzguwGbpNvgz51dWKulWzeyRx2izZlOaMkZEoHH6LkyKNn+T
/BeqqYfEYeOIPBMiopBGTdWrCzn+LKF3tzPQ/zfMRkUEAnsuiTv98Wcn9RrvmvSJkEqB/TOYGF6Z
au00hY1fCY2JzwzF7TiCiJd8TzrMvrI9DguLOewVHD+4AJg5XTM6Yqz8CJwfbk+ZLFMpQH4r3JNO
mHqX0EQBqklvw6IlRSWun9xjUoRbkCj6zVu6SrBvxDbVgxg7ZM+cxTF53YUX/6e0bkAHeCc8bXqO
WHrZm3BRZYsvQ7MJumtWJO6hEauCLEk2wFnL9vlQUZ15yo7HeAj5zW9EHvyKe748hMon2AOhyb4L
ss9edoJxzf4JBI835xPKK4cQAj9wSSRU/6ACbpc51nPNrFq4S5PlURDKRGzvZnLzSyHzig2CX/IB
NHFHQ3o+OClYmCSb5WC610Q/80S/ITmuMf6MK0t3Irl1poJwhMh0+fy4dOEOAcAxeYgELsRr7N8x
H2Ex2NjYHEETX1a9oPjYY53NRdsA6vH91JF4WyUhBeEPGifgx2klBBQ4j8n/Z5QKB3Y/ww5nErXF
S02rb8N9xZ10PBSfgH6fL4kTYU4VCtOI411Jp3mtLQo2QnbXyHLrwDca9s6bUc9FYEGqtJAcVB5i
297phb79lsIjJgUEbGh3AMOoF3wxNZ6iL6m8T2xaH3qGNbcZyD4wzqt++tnVUS3LaaA+Hd/Wol7i
lKVrYt+0pLA0Ucb2a0f5UIx+HiAbsNs75pmtS4Yl8N9WevZI5LQl6AUljF9IOTeIsapMZ8HEgKOB
HrhD5XmpK1F4UPsLqYDxQb4EUcHNIdg6aMLJFZp6MMNg4yzw6gmwiguXcFGeJ/pRWas6wXLFbupa
AYyNWgbcsb3+mrXQJzTuxIqBMQoH3HhnTrC5hZ7xcvtnDUI9J9j4ZTTQiWjx+K4Kr3ULJ/aqJJLr
K6hs9Loc1WtUHRTOfsAFWJJyBCrQUYTvgFxSPEefScxLrBp8uaLw7LrDRXveQCB0bPhNQL6RZjUX
EQisiMmtUlx4To1TBacGWLcl+ZPeqtfgmE1EgDs8AH7aUw4L088xVBXiLqr9fZJzpAxhuQkZukFy
arbUHz3S+QmIpDhLK8PYfOAH+0y9EAGP+oHKDvRPQ3YdAAlbiGj4tLXksNDi3741xms2uPTyvwNv
LGwpobdfryAXQAsH4lx//+ughMNOy30MUBpQyYwM5Dd/fydA75j/mU21+qsIHbosJ5tA3bRULXXZ
T09X4QdbmD+72IPATM+CpSKdyH+BD5sIwa/+AgtMnx8Rp8Dm/MpfMkw2jGP+0j6Lfu2OrdjEJVS9
eYPeeqxOzUZRWdRSI6PX5Xzh/I4NO2qUimejMtaFb349cXV+vvezG+fhQX/DZ38uLxOYYv+Fj/bx
YjEFi1LMD4M0+bSgAF5B/4tCAb7HmqnNOjo9NpbjYfqD33A/k1L+I4/bgafcZRveT3038L+IT/YD
Tij6CMe5WFiAc9EC1dAQn1HZHX9ZnxD/w6KvhBPtBIs8Zy9gGq/2gJ1990whNrWWolR/hyRbJ37w
wmHjia0OfA5ipdBpXa/tpZFhJ4EfBduKUgK1nH6y9KaQ57WWeZgn59S3GAUL7aHkV5WRM0tpbu2q
Q2hQpK2gixGMWy1ZO2KGQeEmoTa0w3iwMpVUvY9aeI7TZv65QV/kkRwgoyb10KYCW0ybvcCBeVK8
HCfIfNH91N8RnGMoAqOdWI8kFF6DVQxSWpvl6aKQMvzm7rlZ+sPz6Gw6/xOvmS4b/FYVNPtBslmh
bM3N1i0ER27ifbaZmmTDMqYNcfIQUT0bJxu80krkOo3Bnz4/c5AKNQT+5CHym/bqaujR+IFkWX+V
dlZ/bqBqapYYLSe/WOlQwdDL7i3m6wgXaCrt3vEg0N5lgmmZAEY72bAV5aN2AaUa9ph8KX4qRl+d
SaWECBHkfmRMuVHDIoPBsMkkbvarNCGCPUxGrNsIYSgDSHJVOGpoevo87OgTP63HluQcuhxxeDGa
CVe9wekFZMmO0CkeKLBshUx8YNZNlhXtsN1Dk2DZjqgbY89AIe2U7HyC6abx8sJWiPTxGXT+acsR
8H39wU71UN7kZuLQTsx8fA341pVVRTZZjisQ/J5u2WsVyFlg4MgGuWPwU9YCaMRAR2CfdCYa95xM
7p5x/bKApDSe8FaNPLepQ3CoFOVtwsXsUujFjZALb/yEjnfAbWrEtWltHyHIqM3xzsle4cUwNK1t
070Aym8st1yKC9zBCS5dEhblJG1tPRVYOOn8ZKyG+xjk4n8h7Qcw4O9mftPcCB3QV0FVWv2/k6MY
B1DRRNC4+Hj/OHL8Ebc1Qt/89101IKvFT6lCeslygQHqmvsCthhZXo0dr2N4d0qztHNvqXtjUI5b
nRyqXCWYFJqRxacS/Dk3vtRfTS9bHCaf1t4fmJB5Ptuu++MFFdNoz6GSr+1MoYZiQ0TXOVzHXFk6
00CXxN4Zu77cRylmB8q3tZkJ1xDYqQD8gQjHvw9EZO5+OCPQlbWgL/a+TkDw9N3ZVhOEQXYH66AJ
kOQquAt3aPiJBufPidzFxP/tlrunm2SbUzzJYP3m1HbWZrijlisPRtWXwJeKkJN+uuIfmdXtVaoT
hgcPUFvXMVF4MTZ1IrgW8g2TsjV2NoGzFrUkOkcJg49DMaqz4EqUyHu/JpfNoZvbDhKc8UODUKt2
FsYyfmW/H1rP+gMOsRQ+ifDrv6tDjYbi/GMQe04SS8JkV4MRDRDi7KLSNx2Yyxhz4mkWueUvUEHC
MfilZERsNzwzWyE2gAE5+Ah/5rFfq97sLbkcDQUeMP6PF0hrr8N3SMdHmnugzNopmcogcNG//nPD
4o2rwzTaL4pbPtTHFJvk4gJbpGIhtGOykzgYnXFMQYaRzr3NH59tRFJKWRzJXFTeD7BNVjvfXa48
P/nnhMDtb6J2C0tOlKu8GUfbqYlmMll0gfnsUFLgpZDzmEtEL8wF1iofKU3efJDa8YNVRsGPtMCw
tMXkq9NiedeSq33WBEXypA+2Shq6G7kN4SdJ3yTUk3sAVMYhRyjhy16gzm+jziVXbqgHE/20HOHd
TBxS4NSC+Ugt5Z4N8cCa6vmvmyGiuK1Vlc/QAQxsqZMUHzaWRPfuB4UPZqCyf4qE/oJIdU6nPTDC
36W/GRCr4MmCpxICbGfnMG9ov34KrBJ3HxiZN+A7V6NRcj+mtgMo56930v02nWaWK86bJMOo9CMf
dzk1spQ5L2FpK79tBMMRnmqO3Ruq9qJP7IIZggbmUsd6a0JOx7tsf9va2fQBXy6rlBLW+p05bzkr
iQ93MtDB0VexmKS6fM4HmU1PEnrL6Qbto+GTj4FEvIGsMtCrB35MwVN3irD4sgos6aEOm1hPBj+W
0QEQtsKC4m6+r74JFcvsqCzP6PSLeGg/q7JeWGazHM09KrfVsdz/xvwFkJMJK9nZDr2LqzHP8Ki0
YVpUDwO1/usSx7kvq3EbaM8XZoiir9IzjUVKeadQ7A413t+CGw3TK54SiPmO12CfHRNTlIqxbsK6
TF/1dVAxqlDVGCslQexda7/VkEeu7lcfqs25sqxk8lNVLsVqGQZvL7U79NZt/jYkUM6BOLCjO3Mq
pdIFb+U9fMcpAKep7SC2h3FKdBt+XYsi2BjGkciwM4z3jCB0+8eHt0SdAU5G2RKfukTuA90g02+5
bhsb0mJ93tvCx4V1bNKu3PPz+g2hma0FJr1Ezv7VS/iI1IjSXQ5tBRzS0EWZEjxFU8GOimqp16+V
aTqcV7y8eQldB5HHiwXrO0MQ+sOu8pd/atpGARgYMdH3wzY/8WCew6pIcky9xmtfRKbRjq1kxtKJ
KZe5QJsOsfQBCusfLgHzMRcAWJaftzmA8tusWHEWGZM6uZiQo50ynBj+8Cb983OAW5H6rcikEz4j
HzENhlGX8exX+uGe/l1xYOdo2WvFFJOyjQXrQWZ1dvtzWtE+i8r/FxDAUDJkMRmfoez4ZlBJ61F+
ucCCLKixEimqcQ0D2A/jjO2+zZwXb2dzIAEtYAzMCZjdAodK3zMcNetoRKUqllAOYLfaGU0ehEcy
SuVlUeBbxf1EUb6kTyTcaQ/hgaAMJqbrp0WUXxoewT6f2gg8prIEJ0dEEq4GDfqRxIaaynintecW
pZf8VI3SI6r38GGF4q9axzso522zMXReNlLYNV6LQJJuam3b++qBPeVw8TucWsGCYyNQk6UjM0gu
lrRp8lj45boFpRxTJmdIyxGVNlgGidV+rfVIWEeylVlMY1+Bb0dPR5nTDSMeKmiDxcbphsu7a1hU
SbsqyE1r+kSX0eatIK0h3iSPuDjWnQ+17+s2toWOIkkciF4czg2i3nldVxHlSDoUq8vNFfG2IKEW
0DG0+YyAhNnkKH6iDrjx+fQoLW2wtILgdq3cSr+fAh7HB7fz4kKPBe6pH5C6fpzNw4IKoT6Wvi8X
+IiCr8aNrzYL9S14getBjTrEBVubKfO/dUUiF0sOoJvj6Fwf/uMwq/kBfG8VGv/Hw3E+mlVnLXL3
muiHep8Pm6nGARtDHAQ5eMeygxi6iEjoPqRncj37ug4kjCsev6fe5xdogIY6ux8D/efttxF71dAE
92AyEhuvWxiTnzZ8xxNqX6NwHkz51q3BE47lcjKmQgQdQxPaZ39687XjRASTFA8fmw5gvJJvRiQw
BIAh+hW3S6WEDXEhcIYvCKWSLnVdKwpbMYJTA5l4x+Ls2e5CR9BknBf1TV9aRfPQxtfqdYoAz+QO
z90u63TSwe3Nkxqwtpm/lKfvG5Yd6bnM0Bql7/coo8r9Ow78tbdEWwRQLGn9OoJ59UJGhsyecXoh
ZuRJCUvu6kZJarYc/T0MeY/llUEfD3NcIFsK5RWHg8GrGEBborCCpId5ER05OudA2LOynj2hNbj7
YDBJ+pTf5hohNTB8BHWaW5lG/6omz4NjQWopZFLrijasXd127jtPyHu2PoThuy+LIyo0kO/PwA3D
ttRcyt926c01GYsHP3PXAw66M5SFoNNO8PIr7UTbyZj/t40WRy1GT7SVWte+wXOKqGzQxkzPD5nf
8CTqZzAvD7Pvdwo7+zR02YPRM7DEQH1L9EHtr8AXYOoB25vFAZ3LmNT/ZJ8idwGSbPv+CkMwplnI
/7tTpXUE/G46SXxE9aDqciNTdrmy8SQXdpuyeSd9rc4HDtaOPXVseCALcR5gW8YXj0CwUwslNxPo
2UWhF3WPUBHyrgfemOIWa0uSNTHSwec8bFdRrSlJxDXhVE5AXg7bDkgSPrAuBy96G+Y+4T4F1Zb8
aTIfcQHL+hdNZcZwpDoagv2RQsn+ds8AENCKZJ+IWGpm5mogYiTMOAGZk3w3/kK4GxzNlUWvckRE
IrQuenxSHN/B9/dXkQNo2wP73WSN4FLb5ueLIvN5s5a7em/XwvOuPcoarxEDrQQkNTANIBY50HjW
sYm6r0ZTHxh0ZqiLB8hjtyG41NwPyz9boOsIFVEkiVsPL9JprTcDvi+RsUHpte3Z6upCJzFX8dAU
EPTQhq1NeiKNy2N5I+wnl6fQL8OOl+adfaoCJvyxZV+E1rUfYIbljP/bOpNfB7jaAtjZvnz8lrqT
A3fJpvj5tOU6gqxvWHdz1lQQeuNFjX90hqlkPEvR3ngsHvsW9VhnqN4arcbxzySJfxAe5tmDFmDo
tiFfBCpmm1ow9mz9q85ZUjIuehAHVhdOW0VESCD1HDCLt696Vkx9+laIPSsjv3g6xvk0Oz56S+TR
C49AX6nkGihzaViQusJK+cijvdlxZKGkcERCT0whx7HAJ8CQLeZaygSJcXo8Cr+P9gZXS+xYqDbO
5MGv5t2Lm+LzMDv9cn7CAl2TfoUeQCeGVn6DhQ/iOvZw7E7mINZ/q8PNAeeixmm4zbkjMQNHOmp0
vmBUQNYDMe2L1bQ+A9YDsR88/ZDFsQ8C3VsoW7M6OF7HoGOJCaT+UwALZs8CVJHhKzqxhUS6GR8J
RCclOUNWCCjfeV2PzC3SPuVZUX6rvwBFzu4QqRyccoIW5DKjgDGaBVNu6O8kKkNu//ZjdYb01CMB
5FwS6E7YAZ8zqL7DFCkDc+LFHaUzE6kHmEIujBEiU/XNCojYwsLH/bZ2OtrpkLSigA42AbTnzFZo
pnBiNgX1BzeVv03n8KJjLXXvMzgKO6sDnrrifGby9NJ2gYdLrj1M7RVbh+IYyFeqzQt0D1O5HuIR
HUnoqYVkH9bqfCHbP8sPKeWL9o7pQYuuSD9j33pWlIH13yIdwBtW5nIxDFrUsqqE+PN2h6mKA3pZ
c7eRmiHJCAlQgLhGss0mEg9fZZ7RLHGSqJShTgMkGLybBLHEqaDLHdflO1YEO5BIgWGWWhlqUH/8
JdOE30PoV5xpQmQlEYWTdur+LPb6vtiJ6aV2+qnXMITamqrIaHNxZGKX7WHQRb3hM15W7Hxdltdn
/aTVuDjtCqU7ZD4pf5otPbOHLhtWkQx6zPDtFbQMUqQ+6GDIgCyD4q15LqjkRVruagMvvidScVN0
D4hYDEYkxjh+ylI5NLeV+EEGfjPNB9LBim5OifrAmTfvKKD6wWUOYl49B6ZaNnsT7L8heemdVD9N
kzIi8zJ7q0YGxhscvcey6tXv1mqJeFXFaEbhO0ENjrrLbJcOrXQIOZIdc69bqwxGvSBDSjmjv4I8
jp36Ms0bgSpwNCB9gPbcByI90m5EDjf1bg3KGwcaqpGI5dhyu6ftJAxponhotqBggaA8Fax64Fum
zxIeFiEFQYuQxrvRd4AgKTNhQRSh2kEt1bIKMZI9y+vYrlRg+MpDHukd02PKumwFoRkri5IIpZp/
uRAb0mUhGQfWRMDPINn3SAiCo3CWlPU9eK4I8RJCGEajnsRAzPzATti/txbsCGOyw55Lyk2qtZWJ
Bae8/SNKuHUsFPYhrztk4+aC/sL3Qci5SPnRCc4pyaLJzn9mFBlcHclsBHpIaKj678JVxXXJJ03b
hQXDG2H6bdQdbCRWGdPEzO9GjsXknKudbvKjLFgphA8ep9Sz/06daS1p+dXHxKyVtEbj9CPMBfIC
0HUN4b4eOY3mhe4vfZ03jpk8BhZ6tX/G1NjQHZU2kfh6Mo/2OXbrCgRDUXnDc3kA/caUr5Iv4cxa
fuTPb9O/BgYwGi4+MJWbdNiUI5zICn1Z2BiDL5/TcETEL2REOxcwHGVSERZf7UGsFNk//V53PN/x
pBeQg5JkynLCkzM47lx1v/77zgehVbnIsmzFse79SW7+4zINoHoULFJaTaKtb3UE426+haoRJ7Yp
ptbEeGkatmAi8UaHtHYPeOmqNzvK5AWoT9vCBbmL/+9+QOvBiCfwCUtQ1Gm0NUhLvmgBiPPySZEk
uUSaitXv6vZn2XOlZDkAb7f7XP2LGFt/g75sVkzNOdD6t1GFX1APBvN9CV2eDTMqFJF32rU8s++5
yNKyAfnMX4o8h9N0vLSGk36Pk6pFYfE5Ld23SfSVNd8OmzJKfkcLl4+qx4+OA4a0PzKSyQIi3dCt
mKsRbdZ/hBAS/+GHvZVqRHxQgI65zscnVAdyRT74p4wTK0vgDtXShhvviOdwuvnUSZFhse6B9I4O
ZBFl09286jwPAIEyKn2u/am88cYkCRfCC7O1XghDRiY8w3CAeZmj2yXuj837fha5CeJ/WOMphyZr
fRFxXCC0PClsz9rxHoNMGCl/Y8StXzmnR9HWGVhWRmCiJpIaJQJRd5k0I6R3LTHSCHjd+rdSv2jQ
QxcF8vNq3kmX1iJa72rQBssFDU6FiswwpZO2o0gxpJCkqn3QX98uKovPGKxeFtdE/mpvXiAGNBFI
0ucUx+NZP3Fcf0DaTVliT3kIHiCHTO/ALoXk1bbyb+tK3gskAi97GeZYJspG8XfJWXJGcZ+oMJu6
LuEb3K2igDtVcVHPjLauxTLe2X0WU8xjDPlTuClsvZws5XBAm2vUCVr2bJKxWd4RW8caQSvjeXEF
6xhKNSNdhF8nEgvAoE/TFOnx387FqujQYgoSaGlEXzLHUdYo1g9Ht4YSeotUCebxNPWemEfPY9Rp
acE0yKB3mX7bsBYuZCPBRazqQQYcL4xou0HBHGPavbhNNRiaRHxiM1DT3/TBAPveMJjFubICtUMC
hwR1zodYYBLwz6mMBRrrBp1sQs0D2zjvB6pnwLiZF0HM+SNEWMPY4R0dxEDEW8sylMUWnIpRRALV
YZvtdWZ0KeXTx71l+bmnfS9Vr7+obyY2WR6AxYYH4KM1/K4YJUDIP5jiTL3MSfRkRae9od5T/wwU
3C/bHpLcYYlOOKiouZSNlElA39hWYKmRB0QAE9KkaUi2gMlbw/5YCjGwQAdqf1zaMPrsUOs0X8/B
LcAWMEntiTi/IiaxBaakur6RfZ1C46a7+/ac9DJJ76wSR636OER4RqDKhdKeYxem9BKFLqDZG6xr
AOoEWjZjryyCGGxh/+0CsMrQTaDJI6Mn6YBY8nXer5BFjyhIdUoHMyuoapyQq2h4WhZpfwLPKyXj
etBbZnBxAjW+2M7xyRfpFHQ5L24wDWAk3ebFsdFiqDIHGqImrKNeZUUAOspTQGq4tSWO/kQIeJwJ
BCK9tsSS3QxCqQAYBtEv6VEzOid4MyWVZVfAaHh6qkYc1mWO1G43ykipGh5XEJ7PtU2MFlngkQGs
ZDyAyUtGcUzvE0tH5IMgBr7I3TdEp/WxBoCq5xN5x/QzMOYHRxddmkJ3vC2X0Y2IJliv4x3ND+0s
UDAPQ6GFGs22IwyISFtxOSbelXCH8aJ7npvzk+ddPiDOIqzFFfKH3fDfk/+HH+XCAw4NoS6+DuF2
25JlZVut/bz1i2hj82remeLOVu3d1jXQ7UWytProEUwZFBgu44hI+VNEew4NvgA4i2UYKq3633mf
wflc6ta+uCmC0qe9lkl3Zathw+6k7IK/KiT2TWclp9/3CrMp1v5iDK8VfeNrHnUR3SXGzCz20LKg
DzndZFK7YW9b2wStIE8h6imjNsNF7egcZsru4tjDqr3P7EcthPN9qg3TefL2gAXBfXCsgt48DdKy
b/RuUHacAQdnZbz/J2V4IZgKDcUiIVCNi1uwtGXUFr7/ao3gbPIcXR58GYFdsh3aFytOuFUDDAx9
MDgJWcixzeQh/LJqd2BACJcSlX7e9RqYG+oYauUFzXmiwW/DZP3gB9pJ4PxNz0yo2pVLBP0dZQV7
iurnGCX7RwmfpmLKKFBqSGZYcPVBIbEIHOxf+21dK+/7H5a0KtsO4dAezLLBsigNENEwsMbl+RlW
3ZioOD7OqGaAxkUX9qFCYe88uRsARs1oxxGjuS0hlmiqpaiZdECcUSo2vh4QhBMJ3s9nI0plvfN+
LoXXEBdBqxr059uojGMjsLMu1gNfbHIYzbS/UWo+eJ5vqCnFhfgFDp12NkwmdlxCJSg2SGhC9kwq
dkIojkHmepWcyTUZKV0WhuD6zJKKe4kTd8Veg+vVOglpXu2LpiZv+nFxPceIdosr2YgTO2agoq+4
FaX5HWR6XY/e8PSSQ0RxQBTaoMS1aMBd13ZjYZQeIjn2YLBu3TcKMugeNaXdL4mLMcxFkN+Ykb28
UMmA4LKIBZvDex4wo9/m7ruA91AeKwjOakzuzAX8ib9eJKz6YvXvM1xgJFtyKTSqGgGIS1FPtZ5R
wtxz5nIIW7FF9aRyHEmAu+kyNipv1REpz7U1tyNHYoVqM2Prbeg05fG7caFwzBHDdtX+0dxDcnKk
Kt/h8ZgtOolcIl3sidE21+05tmLlQpqFWAvEl2O7ZoyqsJNBs7TDNZNoSrhKNKuMJiBxEai1ILdG
wKCk+5l9kvkBbHNH2hnplZWwJjc4ze3eSjgJcKxs3QbQ8XyzMNK0fkqH2GnyOr65otMuIdYUTar5
eXrwHxO9gpa/LaUTLNSuMBKaZi2mcxJbrv2JFbNVar5HzuFF8p4Rj6miOAHMG/jdoG7zOhXxp3YZ
iFT/X1a+gKnl4k7ygh55Ga5nC0+MPcA6WTbcVPE1HScUG/s0lZpKVC9jkphpgzBTTPz6i7Uw4nAb
G+/ogzTH7qcyJNPbZY5gWopoHZ6Q1wW/BuyohZyCBj5qXd/FNVCfS/6qh80XxhuHwGFNbcwrAJFV
4lB8Lrg9kiOj4uagSE+LaRO1GCVxC9+u6JNZRa/AxFshQjiWXu9Co9zxXeO73xrw9a0tkqA5hwRm
b5R9+eQxk9iQchPH9gjGsHTN3Y7Tvym6PbuhLrU4b08RCvuckwCC7dPqm5rNP303GnUaL52SfAvW
vqa5Dr194CP5wRvvc25Rzlk6kuB7lfzQ68AcdoarvVXkVIecrqHsZhfMGdvohHkPQSP3mRUBkYyP
f0wQjLW4wcRco9QmCuoN4Ks7SREOxq7jjh/0zQPLDQ2f6WgE73Fi+75R1C2echp6zyzHuoPavcUm
t9AXSt1IT5oNB6e5uiX5L6sypyc+QooJ8yTpi/OvIKLjudsb1x+AoM2q8R9oR9RoMbSMn9Zw0rhL
+O9uFSNq8EFkNUNj9TnXKf/me4mEm4Uc5qm7mSIuJPL7fZ2/1HmZBG2MG80SzIIyRZSyPp0aiyZ8
6pd+aXQAh4SKhHJBlFqZunQqx9l/cyD/MuQ672bR6vj2nEvpeBB1vEZZwevZCpLK1/VRRU8L1U9J
13A28Lxp5posrDFhCUa18P2SoRpZXgAE1aY56looKfGSkV1hhUxsnPK/MbTvAGFvYpqrmeN6sRjx
ju1VNgMfNGhN1A07GvIzlC6PRmJZ4ctm5QqJRiLe+AnSM+YYSuI3EZJQs/jmmciDhlKZojrYfuI2
QInyH9WAFeoS60gJzXRQp55iWLCGl5qfTv4hjHoC66N3kuz3rstQIcJPKuMRu06pkhzdti/up3BL
nrolF506ZbI2O3MelewQjAdmxM3Y9TPrRU+q/5HZrRN6O6H1oV4dCW9rnUSxM+1rr4FQcMhFPIYA
Wblercpjk8gVWrA0gFsHKWa++TcB2zMvVf+VjJb5TXzinXSHxKD96ULfbrYV45nAw+q0n7za/KNT
YTCMw7fV5FtJn5Xr0/6BP6T1IOdBODAoIkfH+rlUFpPu4Xr07tdW82LlfQNWHgWPTYNY0sBOAHdE
K9SMg8UwSl2jU9NBNm4ID5abHtn0KN3DtDk+BIqeTiLxUazaRCaPq8ffvfoyxduIyz/c5+c4hDEG
x1V4lFE610DsImqgPX4DqtbgQnnPDVDB95O/Hflvjb9DT6QwQLXXOTRaL2n6ffZJfI51A4S8zPcg
Fv3frOECxdcog8z+gr3+kit/9wCXh3CkjzIigMX9QMSULO9MtXj6NifWihyHwcpaZ73e2fLpvnv8
vIBYf1LtNsM9sWd49gtGKXxS3BvK6inBpWCyhUtXBUfoZphvuevxX1RieWlLObCSHFBo91qLEa/5
i/kOR5Gl0Pga3wC8RTl9pgdKCsY6+yp0jTn+7uk+FAdrn0CJPOwWrYoq8bItWV74C4zfCCjWcS2y
WA+WQDd4ZsWjZPT9/kolJYfVncHQx5Y0PdSx6nt3TS5klGodHfIOIlLvKxI4uTTakxGU1T3QNYqB
6VQB3bWhU4lNLJ1nJ72jnm0PFPk7DemmQJZWo/Hjlr6+2W4/t5WWnDyJxRUyVzbf5uhbc6mtiySL
tINZEjvCabTLZ4HquKZZwO8uovpqaNo4qvlNzE/MTv1sf3HUNzmuCOpiWqmbfLODofOjqQHkdXRK
ci5R5L5W9TPtKeBM3nKkJNcsdBWmXlh5pTF6ySUT1JkxNDnE6KFf1lIyNbBijOlrl0yYemJ6uC0V
cAzE4SaRn02M8pIcYZnFsU0YS/smMcOmWVKh6S6h5lq61Wj0fu7mkOvBcPrgpAASYE+rcZZDc0SO
oJlPkGk8BNMZWvUfEg9qhan+tW5GGX0vNZkttpKTKT2NT/As5pkmgkqft9Jh/Mv3h8lw7morqU0e
XTukf5pyx7BtDoP3TLLrQy2unAt2RvshC8+tF43VMmAAuKvxkiPL870xGKRn7A/tU99/Dk+6jL+J
YM0lLnwIww2FWOdP4VTrgnoJiWXQ5lLqTE2UtAxE4bXDHZYNSMsHSSXkLFPzd7wW2PFATnX7k6Kf
xMQxrj9a0DyZjv21R4mDvl/z79p8uag3JVTovHGMZCm5Ml7RSjXSB1LVyqSZaLO6Ek6rJRTc4yJN
9V+TDI0XcOMeWsH7Vmu6W5CwwZ8Sc+C92IDtG8ncF5B1q3f5G1OAr13D/Rq2QHAuFhVnZe4Gl37n
OsDCwLtZx3OfBPnN3SXHbfhzRascUcHe1b1xh5Tz/dOIH1BeoKhP/Aa9AaTTOtvge03I0Pc8rOPE
Wh5gvyESf0bQdV2tWAkQylgFSLx1mIKjaYqPqF30bZQ7qarMOrRlfUXppJkNRFfL3GROatm01fYs
rdA/5qI8c9ZfWP7V962tHoRY99I+7YbIb8iHUxWmytjdlFbMKH4HbFjgPjMrx7gBDD6U9B/vmG5b
LjuFJTz32aVyK5O36pmmL6y6iwg9/wTOu5IFmeJDSsSQ0HuHP4J0WaqhU1wGzL7HIJFv09gzJsp/
9edB+Ia035tUSepY/5XMI5Rh+r5zCRlKNbMfA8q3G6c/fHNwZAEVUucR6vg2GLTXrIbUhXps6Abg
3R26JQhh/FW1Cac2fchuJBeA9EFS6FpT7RLQNEVUtxrUBK56Km5EXwn075Gw1v+ukw/KRdRt+v+j
qlInPG1HKoDFi0QQSwc1p6uNKiuH5GSJmfVv45Mkzy4gBDTZIXLK9ecnwrLkRX1Zbp4shraBwGzn
GEulFLDJnNVr1elXKFS3fEogyIxzVElgWv+ag8R/+dKzBhlD2ig+Ev/AbSWgYl5By4aLyVmVHE7m
y8FZN/u7tY7FgPiA0G7plYMsVNyjJGKRE0VOj5m0SDMteoHFSuWSbs3S3T2TN0lg6mlLptXF42pI
EAtvLTtrfcpEkBLF37oTXGO3E2LL9VsZ4ooKdmO/M5xu45uzCGj7UtN7iTsNnts4Y7lb5ZAtcP9t
TlF2/SKUbm92VLFODTmxa/vjX2RjBl/dJ5DnXt/Kb5/ViAhOhlW7I1fQMBxO13nZ3zAUI2tKSWdl
LFb16Nb+yrjj2hT88fBelTxdothT4ZsIggrZA8z1nbij6iu53t/6Kc0CgYqhWirkN23bhZPqIWE2
7jD/vNKEi/CD2gPncfowX8IgYVTNt5sCGuBDsxyMIDbpAhVTm8qGk9g7e7ZACm6kZ5+swkiQ0aBv
AqxW+bM1NHmcFJrOtwlF3Y0Ff3HAiuInaxIhuGlWkcYbUOCNRqTDMASMgw8vAnZyifqpgJwAbrEz
CpyQHNU2zzP2KFc58RRbenI8SGgO9jtsdltQ6TnCiWX1PHqva/6PDLLqUGB94NKfUYJPpfpfTC0k
C1yf4we6Ss16MzBkPYqKVtqkRJNQ3CgpS3ipJbk4Gg6AU62u2Oopj1fnIMVzi+acByv5MKCFNdH8
tKMGpG2a98BzPLepCN3JQw7Jzbyi2vES+BbySBekyF5UbnWq72H+I0NgKfi7OQXLWi58WMqZkrMJ
Y/VfQgymwamxm3W438Z7mbWdiCgQy8g2ezoxz/yKpl9AL9K8tWBDx7H24BS0c+7cpTsrmS00oSA6
sDDbaTR783B0hfu0IC7up/09EuVhho7ZD4RdN9bT5dY13VyJSXputp0WrPtHvHQeReS0z7nW+Anm
NqtdK7rW9qPF6XQ4Jsf3QY6QUghVvKz+jgra/GfH5uvfMA3sUa+FUodZkechWjPjdUffL3CnKEZh
XlwuaF2WOo9wME2zCl2zN9xbsn9fGkDBvcEq7agg2BnUla5zkJMrCPdimPlDsx4YMvKA9YAMeKUN
Mv1+OV3noJwJDI+r/xsvKclOwYDLXt11TuiDZf1wT7+ab+L5AOD8CZEfK91/uOnWxrUEqiWRzUmE
9tOBqZ9jyoQByn6adI/M2/NxEOl6UPrn52omi8P48hK5/XRHuGIoOremQU9BYx6wiSfdtVKKGB2P
bDbdh70UbGngVxmau2elWW2AM1xA3cF25A2aXIM8ZPOaim0wW9Fw4CwQjQS9TT3wbZkdAOdMC9Xm
aXzQSTICIT8w8zn8nPluv3ay1fU02nvNjLwqduymCJRNZ/1FnOMibnf6AgUmiVPh8N4tx3OoE45J
7vdNNB1ObUOqnxnvMBnhM8G+4u01YuoZRC6IenA9+U4uaZOXlayYDVrDqsjBgtwAbjmRpW8p2wPl
lu8ziPYISGM/+OzJVVqkwcgiBxSi0nFNlQAhHSooLh0Z80fGq2prY6atjDs48OaREzJlXkPtk3L6
LoYbH04P7VV7+uwFnmeN9o276oP1/bXvO9Zey0Qql0I1UaEF4SRDf4PcKmy0t/w5wAoRSxXctu0C
8vnSspwIe9jdhg0So7NsCwhE/3H8x+1eFxZwix2MljMQl60flyxGCtLo8aXvbN17mxcfu/WNB8Lz
xtVFTKZ/DWwhygqb+/3ByhhgNKqwBtaNkmyo4+SlgxHR4gU47oNN8Mkxi/3SQf0IYkMyY8jmB97O
MNcuWkhakc/FrOy4UG1qzU4FiQtFthI73nQsDosyo0suL5vaqxjcA9Igo8M/wtlsRJMC55x1BdNh
jlr1rblaeZp+GaGS5EFD/mHdqy9LYaHRgjp6eU1nUYPgPG3YrcPSOMpShGkKzl1vpckCbn59EwwR
bFXyUPLZ0GI7qD+b1y3iblxhScW1Eekl1JOpLXyEumtkd6tAX1UPpaGeOncWg95U9OmK4MNsZN7v
LT2mBbB8VN+Qiw3Hyb11QsjZmvwKhPqu6ebYpqPZFTEQvia/RRVS7ydI4rmFcKXxqFEEMaIdWoxZ
cD+TH2b7fzPewGyAhBDDdnAQjpYDVfgUEM83Y2x0SaZetufuPKPW51IAf70KjT9Wmxs4ZURmMAnC
hev2XA+bji5JrzbZnYutW8PSh7hC7iRvnUKF1SS7bDKbKyFIYZUQqRsW9uWs00GUPnmUJJ13R1rd
aqCo0Vw+RmevYgdpBxoi4lTR5qc/yLQrnTgq5j6w3oK5ik88Ut5apLcSKqAwD5Rzyw/MKV1wkdVP
j+FKcgsCqZ289JuTCIScaKCbhfig+hC2kmeJECS0gdNNSuLBJGDoBwNh2DyGXjBP4YKzeeQwKGxV
ykBIoU/kZPfu83Nric8JM/0rnqZ/+XYP9UQuP7+ul2in87twgWm5eKXca1mbI+XLCZaOAtFT75R+
ApsUrHEwRlKeKD4SGnhdlYwTkqKLXQ5FdnXwxho8ZZhOAfv3cHKqM2YPVbyeaLGrjDJRGI1Uju7W
b22qCHcIuHUhXj+ZuE7hdeqskTUxinWwNHwsaxjBindh3z43CAgmUGX3X5UEuPCnElpageQx7Oz6
T+lg+O1iCjCpRWgnLqhKCZuPdVBZeq13upCT/ZzIsf+K/l28NQNYTZukn6Opb1yFSsrZNGzr6SSH
/THUkrLkIaiTyA99nVprcPlHxiWR5IWXb128oTyXMcP0ckYpgFthLH1XAc09SlfQOf6TB4Z/Zmu0
V87gk3vjIEbtDJL/sjVDgancffyZxgqCU+EgN+LfuL+KjxblBqEFXpXawM4E6wkbArFA5Ne/Azeg
D4Cw0mu1IDtkz13fx4njOHsh6uFqgWpZxZcC/GF5dW355PvfNKZQsVKb71lPF8vtOuYObhy4uYXZ
blVW7cZhZlKgRPwak6SPlXqphFo2bVTbUaJD3Fj2B5r+r2pN3z/kPIJHe/2wzwe1SPQemw5o+Lor
nk0CoxyYimLv45ojw8j45n2u/3dAe+o9lCEnOnXrmhI/20HGYvUddfUmx2o9J3/ENgHksqve88Au
X2B++XpZ9RiNeQWP6ZnoBBxe1E5z4d5iOkuLSLVKJ6KP1+RQ4AhyRDVQs3hMpgyQoskid0O671YE
nW+uBghWuMuEVxN56RG1G9hfh7VRz2lgB+6rUOixn87MxyQWWA2sL9wVhJSKxShysK+BmSCzubfI
UMFYfyEk/r1Jtug+h0YGLlYhegVcCilb5SOUmgjbxeo8wQsK+u8P3WfOrfpAA79TKV/icOKgHz4J
LBQ5quC0SUiSWgEz9RyGyhdBlEgDedxXjZhnLAISQxkPi0DBxfAoCwjVPmnAJKRtRWnM7kmua9pF
dIlUYcPkLNUIz6fFC4o3LX6UR2/naKv/8hL7EHxDB1e6TTu3t9WMaVU2KrcucTX7H8l0pWS7P/3s
NT49tTEeptK2jFmWFF79+6Ig+2p1t/MRjIL36sfSv6X+76JAarGjbaoo7cTqw5L9Ljlnu4jjUaPz
xBogAM9b5bQVS7mOwITOotM/36tzq2B2POcsMsyVmhzOyLuhdQqt/TQT50KwCLJPGMqI+Ft3cY6r
DA38TQ4cpr+rypr6EnarqYaTGW+WpXpOcTf4qvA7kXtsTOc3oMDynZk65eaKz1NhxEBhQBEmbZFR
eehT5bnccI37/MGExJSkzR2uFRvIJgXKGVVPSJZdcZDNBIL+jVWTFNj0x9ego9xWC9VE5K/uk1TT
KyHehN0O1iUQE+2I6Tkboc7Y7VYr/3UInz48jorTR5pO4Gf9bZoq79HEBqWGxmgUHyRDCyg+eoY3
gmZNI56aSprRE/ZbQBVLDHvhCfRrFg7vV3Blj96RGvVRjMrENr8tjTCATv3CMVUI81btX3UoJVJa
0BtunMaikJv18uBQIzCagovtTb1aeSXwSssIerLrvPeqZVQZk0nJBqx8TPFG3p1kWbJM1a9Qlpee
tlkuXKSIXkMB+9szOIXvm4m8u6zYCo1ITal4E0JDnRTQ6FJgZ/i5SZsHP8IrUM7a1PHzeM7fmn2u
uZulO7MfUYw6Bwqpm7q9hQF7BJQn/xUNr12uhVKVvatHQpUhNX8oTT+09rnspGc+2RR7A4LKdUk+
0xcHqrYAbczc87q2rfcsmqh4RpBoa0UhuKAjCcYAPnioGO2jxVJBZXPNz/y/vMZTfl4Nv7V1hC+i
1h9jYRzuq5OKXJ6wHiycPZY1MMVShecODN0MdR0k9NiK/er0P/5zK2MxvD2Bj4WxvOYJKVZouqK1
RT5DVH6JwyzcmMLFTHGVbzLQADKImhf+ODj0D4wnPKDl1cMtOm5y1eYKGTy5KXqxgdoGh87YAl5B
xiQME1FfBJLu3Bitd0EmpQussdvOY2OCwitCVhrjs0CzXlzsdGCCpTkRs/05Bp49JYXb4P+BmIC9
bvm96eqoXAEWe6/8mF9x4aHi0M69FwuUHFlLheDsKmPqaeB3hosrooq1B5obmGlXIHVT1GP/fJpT
xWgnymhCGlL5rcvxLf64RKosYd3Ub41/GkyXykyUk4hPdplhRqSPCcEuCmdIpw9/2K9kgR6JFAwh
ITViNFu/SyBfjOVLW7PGtYbA43wtJB/5+94jBTrC6QJp/8xJaAb8vzPBTKBUahjqqDSR6gH4+3Lb
aeScdffsfVaU7tTfIjAcCaXLk4wQ85EgMIROPmWht1dVX7lCS2Yq4kDCGqlsddA0mdLNtnpSlN+J
4FpXO6meX025oEkG5FULmdYlTL2Xpe8rkd5w1cyrmmfe3VoKIyXc5qOUMz8N7NM9EYVYJB/YwT1G
DgJHA3vsqtY+KpcD68Pasji2SdsDRFKzHbSFwBraLthsM2oYU1bfM5bNhaVGndn45loZ+DPDJGmp
Z7tKi1jGPbBv2QYz5P/CvsFGYytaF3fojSwHUSoT3RX2HrYgykZgf343QZCM8M77V125xallthJw
lBtDApFp/ka8f3TRMUba5tnYqARfUnssmNA0mLoYxm4bJbTT2D4fvjlvWqr30XmXBsd9uYUeU9jk
JD+gGypzqcxNLXNlSNqY0jyPrgrrBJQDd/T0DRAGLH2OjlMdPodivEb217NvOcaMGNIz4EwlWy86
YExFYq4MfqMJjdJzrtkEmsaTNnGM2y6i4N57lELo2vp5aXQPdq5yMI+RlqBmMv7pb7k4VE36n9ib
i8cF5w0z6knWmuXG9lFR/mCgEASVU9jy2WlvcKp17XHiYOGobpmsPnPr92cOAYX4XergZGVNRFgJ
H/2+I3B1Ajf6IxDKxvudgl4WgFvszQ4SGLecWpPuyL/lwO8+fh+KEFIKzneX+QftIaqaoojhqHHF
DHHzUSui8dMraC5Nqaeeq984/zSMzS6EqUfbhSTqmZ9YeY4sJTlSLIv8z0K1GTU+gM9DDQNOnIwm
IgGIDzAFufRLGLe9LBG7XzlxPiTpXpu+aOyCnbdkU83MpjL8FrbCfqkq2fkKyOOcFl+8Vct6/koN
fRWbAlpTon+JPE2wV3fKdECVeFNh/iKyZE4HNMxmPvf9/m+I2ZcJircJInJTau4bR/Put9TAIGZJ
LPs6YVi8DXepQXgA52ag2wIyhPGTXeK6nXUD1CetfGMBzhWPkgLzYyQS2PCtkHUkwyTaMW0ZtaC3
Y+MkvO0I/R0KiDt9FQS5bmGF0wI3AJDl76TB42rqDa9aYmVb8P09s8oi17XdI7gg6yeP+7bo5BZa
osEQ2lOduLUtwh+DFiQQFVvE3wkfn1N1PfAc+avcBSOj5fFOZapn+9pG4mYHBpOt8l5a8wjHv2La
kPVGracJAjBs4+BI44IMZaDbseZp1xBcmX4p6J8C7GtxWBmUl3IZPanK6DWPWQBShjsPm6RhfI2g
zUsIzkOEZZLfMMaoFI9VDX0U+x/u2ovpixlAlEE6ywllyEEiJBOB2nWMKxAZWyGCTGtEk5Kn5w2Y
WW16XC6mtw0bG7y6oCHtEx/iF+qWsnLUTRfrkrSpBtal8PK+VzhScADMSaltk+zjzkGMGqUGUTW/
UX82cQjymSn5ApsQQD2nLndC+jZoW/pQJzvLCjFx3NS4/I8NuN8e6aHUeOqVyERWOoW7KL1FRSjw
KWDUeT7ApqnS6Xfqaj4dp4ZZSl3Y6XdVWDpmM61ysGOHPTgkXsDb1xYBDcjZz0lgrDxyYaJRR3Xg
OGb5XAk51cpQ8GdjPE45XA0aj93WLGstACpni8VCCbZm3sobWjOYI2jC+68daMsIUgzPWG79VgAj
Rv8ZPAsThjDiyFxqK95rS8NSuzqnAmCJUF8yK+MM+amUVWYVq/e7myRr+fQPoD4jQorvGKjhZKFD
uuj3pBVaPBoP/uyPdeM33Tg4dWvPYQSSz0uY8SmLO//qKMhPFrLupHRWsGHOrOd1CLM8KQERND6b
x2EmAyZvvtZXmvAGsHMAO+yerei8Kfu0kU4rCohKQNIARJJwncjDnBx9GPBUEa74F4pn6HUP/kQh
8ff1gpmNP+QHPbEpN6YIkBq+UD2NsWjoIaHuqMYzGezVsoKiypZMGfrLWBFqPUCCL6AnEqtHzLSR
F6Tjri8WQ6mHS4WA2vTtZ1QwW4JJxR7t4FUKANxHvOChLoTEWZy5hGwAxnXRCi6BZhR829ktlZOU
f4+B/WOxcVvmYFbJRECr9OOLstpFBMN1KNSL1PLBS/7B6ZMk/8y22prUYGfQuksJXU75CTzTJzG9
kHXwzO+Hb6U8JtVlvhmRUdqJEPEyoRt9pjtIGpQL4K/LHXLMKS8NEzdLsoBm7ZlGm6VVNc1fnMmH
+2Go59C85qwLXl0s8n3LjYnxtpIoO5HQiGDhs2te+s6rjXZcV+KdeTylTeeHrQpVjtbvcFwJiEWW
vGrllml6SOvpiTJ+KvtDQZDXMPdyK1405NvgVadEqwymuumUFZdke2uD/aztemznw3niMDLRsvoC
/6STBzn0xZ7nb98QJ2PM3MApfb0ZsCNAskYj+/4iLIBqgcbkBnlksfDBdt8rHKScfMO6Fh+aV292
SGhDDf9GraU0HweScdM9sJHmXAyBmxxpVNH5LdcVqBp3Zthi853CqHmzb7mZLSzddYnwjMarGuti
5WvvyJC6IBGoGodOXCrRSN42UkxgXfSUSn6zX9si6vP8kfuHKbPFx4RmlhLfHryH3Za/hTu2PU2r
0y5kvhDorxtpYSvC7jcaX86I/D1D13Ll9gOYN60od81hxoesOUVLyh76vAqsu+xIetrua7rgfAGA
7djt4dbNHObgpf0MGgmYjHlzCFOi3YSJ8JwL3p/bL7uOiTfiyncuyUCaELHpKUDCpZ9DuZNq44/d
URUNXj3qNNTFyXz6dM7yUiZiqblpollu+T8b8CEI4lHI72YL0koQhco6MlRxs8gBVF89/ng4j/7p
3hUodJLFY7VZnBH/hMSvSraYDave4Zzhlu0l5ofrQDkkqgHIDpEpyHUIP4AusN78ZHpS2QeWU9pf
W8ERNBTLY2x4hL59XVhQ4H/V2E5MJICs+CZV9I5YBiyjI5Zjy3ju4H8737xE7O9qYC6ek3Ccsb0q
w2mHCsCfzqcd0GV3TErzVmH64Kgec5VJjs44Hq6eMobKT5/9C+Ilt1Fg8pqfGN2tgpSi40NOTmKS
U3E3ihqnTqFA6coff16WRqbAqn9p2uXh9kXqmXaIFlUjW/0lvnWu5PYDv4ot3oGVI3lD/aURqgsx
GBb5vcVOUic7GLyVNB7xRipveNgpIY46qlsJchhEjAowLbe58IyEo1Fe222qqpMjGpS0S/UhL6Ou
bOnjTbpFyY+wrmAAy5Pwk+STDZSBhqZ3q32zzcJbVq4iiTlkKJFTdgkkBbnDtrayRgMXupBfl+Qm
4re2ZXKLLQWJg2rrF+GsSJfRFDJ/eVGedvNnfwuj8MsG/2bvsMnfa1qSsXIXXd8rnu6Z56U6hNwk
i1cLGLghHUHmOtBmbBkWXkXEBc7st5KgYCIr1MBXecSs0Ij/vMQDseNmjAs7VuSvvtfmJ5BEN1Co
Ly8K/UaJlhTUFOOyGPD8UWzztl2gTu1pYPA4b9w0Y5cAvYp0/zKB61ZF2D9uD8jWJolrLNAESmMP
A+I0evQclM2NlEpHsVCQlbUeaPkGzn25eFtTYLNmBfRkQJkM69wUbs4rvpsJYsVndTnaTYmTbsx9
vcI36k22Qm6SVXNwOId4Sbro9ZJhRoc6GJnVhHlwKS/VOuVFohuKeEJUrbMdY+MulUhIDdPXDVqq
8Phkso3qo8hjET1l6OBxRYpr/LVFcCFobpq0b2qEpgH7E7nYi3qA4RHcIiwMU+vBeyoalvjrUhG9
/uGy8j3g2JDhHNmIFR3T0EdD8841etkH/bnhMhWhuUBulcXp1wbyWwPPcGioTP9AY4dMyeHxwyEB
FBVBcfYlRZ3TkjNo5cVQWAyNvoyZnHqoo1sR024FY4zsibuWsrrQgm0luQ5B86y7syBLnlnmTFkV
U06uu5JU2Bm1AHffr4bnd92yV2uNj2Pd1c2QIqUSdGCAhT5n5IQVh4QxojSzpMubrX5udStRkXZV
EKy2qDSyweKfWZk1prELvyYiqV5RlEqxJOBhJ/LXJ0dCp3zpVx0LGPnZmV2WlKJI3Dkeh8QDCSmY
M7meU4VuWTPoguZ7mucqGZCRtG58wtvfp2YEaqHc14wN1BqRvhRQVQ7/DD4mX+/ZLwQ2QCQoiCfU
BFHPQLPSIg01Hs7O4YIi92awpQX2gTuFoEDjVEKppHad1f6tqb7Ep4bTA+D2lLuIBvBay926JUOU
bz/7GNyJv1K4apg6P0zNpBSVx7Ecb+7KFn0N4tDoq5O2Mi30gjUmFCWSCMfSiKZ65USk96QAYsIH
uzvS7uL/56NdEDucjpOkdDdorhpWcUH1M3Kc2zFTd/SNYwh3hmc5sr9TXc6ecEJfXf3/cBi7+oCP
JiuiGQFLuriwko/OUCDHSZGbkwVQXGJmj4acC0E3ap/jdWSEdwreTWONDdsKm+n8asXjOzEfvvlM
rJ++40N9HG+sruKejeVGVrqSBPW3aGH8+eHBv0zCpWMQF7x+CMYCwElwPVSt9U+i/XQSmgcyp7nB
tI7f84cRqXWO3+zmisO+TBluyn3V7rtG2MzNXne5pCr5l3W5l80vwPsCiDr9asxH9GPTM4VGm2yX
akdpy3jlXNqsLRSvYAqA+21dTSicCZwM44Pai1PfmuCYKYCL1JWyqEO48LGnRdAPgytYBgQUyNec
qWfKC2sAk1z3SSAkvA+tBJUPmbKz2kWjYycriUgSkhWj/1TOniOsHGCAc/umw1mZmzV5LAtjEoqj
dZHaNy8oLn1PBQG5OoHOoov34RXoJU9kR7sOfjuWiFIUEFKzYhwSBhvwGPwHWvUPFtC2gGUsn89p
DFeQfZgIFLdsS45jdiVEohJYQsfZRMtR2E7u9/wMFDD5HveMIFT9dJWYPjW+NAPsP4u16RlgWjjN
dcM8jyHV74TMrWC49tCSkSDtlB9hTO6UqhQcMu2FUjlNFBAgPftkz7sDQAE6tjC1B5GXGmpu1oeK
Gx8DCzS1AmQCIvrA8StWxM1pUwibZBdkulMH6TvDfpY08pegkCHfhoK2mQArjpuZwZiABSjvhiIO
IzicUOVRpM5SJoZ5I1qnRDEwSiWzMO0FltKuk/jSN55afiaU50bwRrAc3FgmnEolSb7HhB49OtuO
ShHtd9vSHwh8ZpqwFGlRTIRt9cYzPer/3nfmBcTGGSCwi2sYx4iLuf6mfwsd8YIaZi/qrcn8o4Ik
Yq6NB/1Q4EcV1u5vHWi84/mDeJe8B2wQeT4l1c/LfAZ0N7m5FDth3dRrAhUw/8AOG2Xm7eFfc5vJ
9HttwcW4FplZP5lXbLRUHEn3bdpSvKeTB10mT23f3zMJhyVJiXr0GPwq4N/a9rVcPyPFUUX+tU/i
Vw1wxw/5rDsd74OheasD3sw/NjIN1KZnU4cCCSiyRsdOLTibNfoBQEc5AfmuKJWKzkvO8Dm4rDoS
RvErHQKi0rxqo3MtvLPJoxsCjIU8mTN9sqT9p1Vbts4ADo+8ogzEEw23kxe5PUPTCe1cfKtVdrdh
9/ZDCC6nM7a7dNNwYoIncdXae/PjiqaoRr1AIplZKNsQNeHa/jCcS04zaMn0aTJTJ2KeVZ3s6zwZ
/1QFmrblvwa/wU0LtaG9ZvVGxfOG1RjXAQmRtPeBSqIFOEXHI9K94Kmo7oxyDw1SX+oUBj0v3ABq
3+COvd8JPGXLoISWCS4mk+O/qZWoP4GMxfvVR97rVrULcCAWe3+nu7GjjC9U0lClhYJ8DUkmQB7f
/McKdwsoqJIM4VDFb/kYAV8Jj9ROEWchbSKJURGa9eW4zHK9wNBMWvW0uA29S4BzMUnoFgG9WPV8
TZEkR/Y9CbEXeJJYGQwBg5cNq7az26D6tB3GGgYa3Y9yozLgHW5I1BvxHSQTbANlZTZzRn/W9TSj
ieiEgo0sTcHKtua3egxMBKxyUxLSbiLDDddBVFWKO7XtX/JNXex0QwiGd5+LHxQwLCqGOdo9dUSj
r0STLmMjlQ+Gi9F0ytZCRl0K8+S28dTs3iuVSdykjz5vEx4zvIssv4yI/QaiilN+Vzquy+Qq5QBS
FLWmjVScVovNy7SjGeGni61dZAWnGxXyYEKj5a7fKr7NlI4VdxS6GUTcLaA9pkE1iBayOQs9BFIF
ZhnjHYPclQqrDgRap5oaLx+rYWEes7uwwkXiZ7qwS6UC73abzrpnLyIG3hf4NU0AYJAfbP8rqRGe
VTeCtkxD2j56LRaQ0EpvWzyE8CGR2mqQP82j4pvUHooOaJ5moIRqpsVT9ABBgSm2GodlIkNWEePK
pmt+FkkQnVk/BBnL7v3uba4S8Ypu8QPBcRvSbh8L9IbYcpT+OGYzt+9kwjo4qjlEcUXeQHDzPeyG
WJQLwnyY/bVYHBAHjupn8Mtyznx8RShHQgqshV11xGzUq4XzZtjR+dUnz0St/OLVCbuXXWnkgWNo
g6rnuoOffuC0mHbf1EbG+iYb7xQihb/mnHxuT7q64eWOBxdBnsB1zHFkgwRdWNJt1tqeEORSqBwA
kKrQYiEroK91HppWSDy0Pp13l8hDdtWnH/Qn0s3kkuLBuleP1vtZaoeVWLJbH53fAQa7nRWzf5yt
x9aeb56z1GWRmsQCVt+LqfWG3MoWzTmrOAlG9zeADYeps0iWN2/w8l4ae0jK9pz8o7ZzDDehqVhq
y/7FUOUz+orNO9yTI86fIx8Gcoq6RzX74zXiJZNbT/O/lSzYg8pPMz1PSkKDTsQs7v6zXcLL4cIA
9jRDtEkSAkzm/tXHVHLGgyrZfpfJbEQc4ZFC85Pvnc5O5MVVko3fJ9Sery6lg6d6HHo2HEkD2+AT
iMyQbacyA4o3peajLpD15OyNuAx1mc9nIDl5aqUVxWS04310fx4SW8nMvYPKqQ3s1nm8e90Iuj5B
I3rdPioJieYGe3AJHt4bgHCrsrH8UQFqEpS3Q/yRYCVJqidLBASyKi7PLAzOtcVOQOS5tJC4NT5a
KeHb/cppdD2UdOQRV9QkenOEwo0BGdRvOEQu45cZfatF2NsSd0KFfUtiUMrqo8WLaQRCQmJ56NFG
3EzLZY21jQk2uqIZVXyQ9xZj3XltRxhFcSySR42oo4jsl7wiN6zBH+YoVvG2ql+5BCmKpUp1XneJ
k7qxr84zT2nekWCRKCM6JSSshyIuH+pYIfs6J5hCGY4OJMQ7vuEPEkvvVK/RB9DJ666Y9uNBhszf
r67Pa+dbmr4I3X4yF8n1vJZwJTRhw8lYtrYrlhbeE04NzvKfESNpr9+Y0yTJxRdR6xNrbZp9q4G8
H0Fmlysgp9QOaHjvDI4NPInDfJ8Emq6vgQTBS8nEAAX7pS76T0l092AQwjQ50Wj+/UISoAaOeGoR
6yW7bwFfd4Vom6LXAcGnlm/P950/Da/EEgrJBe8txRgS/HCSZxNisg8ljidByPeKsWB3K1JXGvt1
PwgCOdv8OKqCemQ9QecCqmndT0F+G9cApge0QpBxQplx1xcx0ws1gZ51rHTUpetANbgGsfJqJxWv
1Y22B/si4V5gb9NoyUntJSDLoO8vTC1hMPawRh9BAfYu39bgN5Iw6n48lA8bqABTS77Qwb1KDOVy
NPwzQRFXkncrTdh7YQ0fh8i0bfzDaTG5S1MOyYy9qEQgSoFJ0KDesMC2/DmbpMwywvl7G0QhkGmw
Bz8pKOsYFy72HAlgPua+SNzc9fzlDAfl4IVTD5k5cUJsboA93IIKVNX70baalE6Fh435vrypwl7v
hzf3dgm6rQ2KkpIvVMF+eW3i50gqjVJiv08ztVw2JcB9Tnfodpz0o1ub4l/+STjs8dAVY2APbCwp
jjbcsS6rdJkFgGlnn3Y3keljJ2NIQrUS0PWmtHDY9P9zVKef7IEuW7biAtJswXUYZ7RJ5/wMKKCr
NY1NTaA43/Mjhp1P1uvzeArFihWeyam6RrQnFlXRmRZvvQDXsADBVPpHFyIvUYQBNRtRW86YzPSy
WRgFuCWqiqxWVTW86L/DTCRqwHuE3ZuOvqTXL6y5Er3sYiHCdcnsroSoC4YZ/7mIo0tkJHhvJ2KD
HFgX/HUEET1/UaSxSBzB6Gm0Osg9vsWuBPosC2OmsWvdmw/4O042CDLnRxqXMuiGZPZiB9aGUUrD
ozRyQUrgyxqnHRbe/+3MluKhu9Yedv9YODpY0A7qQDCwRhVyTX6TEwxMQnK5ct9DvWUnWvCGBnpw
+EoiPhCgawIa07zPu+AC7kXjLdvi1VoG939cr7O00cxuYmtQtrJBoKGf88iL9I79pXiOAX8OEHRX
hH9e4UReA1UYEKKzTQYfGdgjYMC4zRNASxQaCx/HDGIyVOCuo7Xb5Y2KifsNKn3q8tlg4myex9Yl
/78l6P5bYS5zFWA5N0KlXv5Pf/6M1N7VS8xlL52evvO9JoWajtuypE5Jhr8++nnD2pj0iH7+JmdJ
KB7X+7IHcoO2KMORe5zLx6qih4ALkPHuXKZoEp5lY+SrYXwRLOvDK+yK7EB0xQB9bY983UXC1wRr
btciFT7jmdqQ3GtvFrlcmsBEhrPFr5qtzhMHlEcnPzqnxJwmxYred1WAPc8vx2y6xaidxDwjRrTt
Iaz161Ya9JCt4cKcn1WFefv5m5H/INdiqM5IJKw695+ywBvSOu57kBTItNxFram80rbp9TaARIgK
gfbDsWg8IfviG4kuccmVgmWFFz6qi5DIWY+qYSjnzyIgJ13hiST7RAwxcVUGk79qBnBrxCSrgwL/
7q8ycUGWoCOzI9QSooSnw1bSTJV3gwhd4npkeLnchy+D0xKK/l8PsLd2mIifIuiX9oxsbqaN5kfd
dvq9nFHa28YsHQLBKxkVQpP6ag4n5wPvwlkFv1ERBknHYRK2VorrQEXR3GUBhMqe4i3rHFq8PW3/
dtiqFpA2Nzb2hEoEjcyIYftga4D+I4IUGro75noiyz3ktxRb9pZI3uZyUVcmKrIkyJiLdpZuQ8qM
Fn+jSc9zkLmfST6XQigsrUmxsJ2x/h9hI0ysVkhKQRYufBVuBcqz8bL172tsRBWI1HX49ctBiwHh
AvBu69gJ+ZsIrTTjMKkkm9lFEy3R/2wbW87ISU1O298gP8FPVftqUUBKVepc03Tx2nY0+I+Jff9p
M40vaZwqKT4VJP51sEfzIdrokAvM6i0+4YVAQctLZSLVeTX8WYk/0yIeaBjfPCLnMh9d2Hc5gttU
2xCrwqhHXuRbQuE4frpjVbQL6iMXTl49p9VKoKRN/j52Loqv1uV9Q4X2eJiE8frx+Ok5qbKo7Gw3
NoINJaYqIa85Ca4I8Pk+7tNCqmhunk4+32JOKEvIpUmWRR+bJwz4Nx1GB/NxgCiQPo8pVNijbMgc
fwUriAOfuRHXYh9Vb7X5EV1vTqfrnHBhTjVlMwc0yHIWnq45XJ3XAvHs9XVWTlU3V9o+sX3cs9u4
3A/xq9Sio5GPXY53PPLbt6cSm36+8KV3RUpFgNvInXKVfkZhDSyFS2phTKB4tuV0i8D9ngwqb8FB
dDHbvJxZ/92n+6xFVTbOIoynGjJqF+6fCTOWixTUjiF/s9bXcIEOooFgQ0kLVNwu/AX0tUZjLGkL
a8h7wR0+IS6qQ+c2pQQV/tkElMGKA49QC99AZL0WDn1Cz9Ey4CtqGDsgXgdIPBW0B5Jbg81swqSi
BXgxVT1R0K/nMbXRfcW4lz45X+s48y4ePZQ99fr7CYm2iO8T/XVHr9NxCPmUqcjpaircYiRGgozx
u/ipSaqb/Rqx1RM5xNDsHIbTYFzPssJgAfis2TJkCQQ+u1XabUAimSIO+zxZDlJWi5BraVLFgQlQ
+/XEHH7/9tDsJ8WN2trGvfH/6QfDV65zRmRkBT4rLwQdU+1OArwvTvF0/36zQP7QkL8ty0fjbMOp
51213DbjIP4ggOhHCumYwFJIpSoDX1XZaMVDQsdNEzhrEmLFHV6mZl34p+zIDnkQ5tLauAJPm7/O
PtRxd91ilBRqr/Atn4KXhON6hC30nogRokfSq4Ka53D2F4TCdjhRjzlIx+X4W/tfIYM6+j5Xyic6
qcQ0mwOQR8PjoM8Xdy8Qn4+EUVPGZGdrzIiiJkMs5w4CkTg0VXezW2LnCV9uj58P8Y1Nvm9a8CoF
BqMTRWEfcQTKHN4zMmsSBdNVAusuyK7bGSK6OZZec+CQTMbUFJlBXo3jOmzlrJ2tKE11a96n8oCV
gZqOykBjwcCeqsy+4KHpkh8ELKEPGjP5oQazXFtHW50Am2jG/hYs6Sh0vMOFXOmVDMFDPeAbCzrc
4A8we7Ix1dwcy66wTrCjIUQCYBP+ZgpsWfsFDD+lOdO7T4jXxsYSr/vLjrN5/4+kKm3H8/GbuYmH
iwPDLIbetz26jGh+4yZmcT+nzt8o06fd6kYf4pZZRU38++UKPtAbcWosvrutSnTdeM3pov/IA/LN
Xr4fcoFiYeQP7PXJP90aaxEhCXP3cy0wjDbPzkIAY3oQBVhxxoBaJD3BJCGtSBqowEWLezaBecea
7e6+VO3v5bJh+RzvVXbmob2ecyAAFz84xBItJzE8CAIBvSwLtlHv2aos92vHbRuAml0U7Ge595jT
62v30l67AsfmeeHfWjM1BF3+m+wR4lfFtZYV0hCIdRTIrf7Q35T60/GcCqEEyFVnXd5ddR7UQ48q
9M0M0relvhWx3ssG9i5u/GRbfwHJ4DV2go3Y6NjfRQACb4lJtnGHCn+aC8Y/0piTpNV6nflG/iem
lTokurBV8sqVtt1srltYqVbXywvtjBsTzQC7LsKVS9qYeua3k8rxl3yBFRlbbw+QtV8JgEFlxSLE
Xdc197DrTOOsiVrUiiQGgQUagyaCpkRgKWqPCefQNSgMsfV18aexR9axE5cqHqu57TZ5oncXLBjV
C/nspGLBg0ynZ4S9euIOCDQW4/C37GzXX1+NcjShdLvB1QOciQ4FT7qNR5AcGRbNOJw1dHMjFRzp
Qh42keGeDGLZw29EhYBkX4UuAvsfBqjXTloZ/Z8PTvUPRqltN89Gd5ipwjsts1ZzT711/RtZaz+U
i9+t0mBeiaiXFAzCFuIKohdpRQbVWZODaDJlCY2f6r987Xhbqxx5guWP+S6/fj8FbxXnymnkUXea
mHgLK2SFxCSdNZ77+o7OMTwy9XTQvN72csTir9ejFEA6yDWZ4JRU247rCU1gG1exJ+Awj/FcVIRQ
DGyHiLaYcPTtmDS5Yosld3He2tShODvGlxjNkAggntMuz5mq1ELjHevgE4Eje0otXwCwCko8UgiN
0c8oNRwzyHkWX09tOQ9Z+eGIFcG7NIeq4cV/7mhIV57kC/pIMwWRB+oUzo0fKwHHP4fSB+X6Ko5y
ITmxStohA0S8Q1/Z+wbp0FQQHgkNivfu7898BEJ11qp7+F7ACRqdAHT5PNxIcVsmSb1eWXfmyxSr
nUUJfua2noAGHRGMbWTJ+FlN8dAYE2iPM1XGyzfSF/lns1f66b0QFsAIl01rXDbE1mI5HlhKzfn2
SAJE/8J3cA8AT2FY+BxAjT6axhWdmiTReraa0dBdMNz7Rhq3M6W9lGKxc8LgsHZ0E0eWxgg5fwKb
ukfPvVyAKAh+XZsKj8iTOvY4oKzSm1SPp4Bkp9VVcAA7UdWYtt8fzZS8NrNSEg2/3FrzbecfXl+L
NghqRsWztfboieZ9B2MFJIxq45qdnxsLHQ6NSOCKU3nY+P4cVaMc2tBsD3S8WkOot0OWkn2bXA82
qz+Cu3J+Z7HKl71uuKRJTIfV4F58LpiIjZVfIyXunc5qx5F3BnIgRmT6TluAKZzIZxSMPRoFrm4E
cNovkT5a+qlHGdrot048C9glwDnjddAdB1RiR10E3xb9BJRC5fU6PRvtksS+gGfev+ymbKncj4jS
RItWFResSE3TsKhinB/pjjwT/Vns19RE59uAtgC6dE8kJKqRgCYsdXvctbe43dg6H229m6/+e5qa
cpD3z93sB1N8fsllOHc2Tz5GlANJ9hCMneDsO8luf5X18yjt3mvKXSd6a0qCsKY2/+6x50e5JEO9
EHHFCmiZiY4WFd5Yuu2Wpp6c93+arpma9e+tTLWgOSAnnvp0QW7zRy2BTvKdt9u1Q3mn6EziIfTK
PMnLhTNwD1MopOiW4rI2A6/tfWKzcqYTMAaqWuRJ2/M/LbUYBTM5E/falOsecjaGWo6WESXR3lMp
Op3nOclD/H/Xn1oliKk7L6GRf7KVqFJ1yEGrmkZxljTuWiw4LSa6fizTlkRtwhRPaQhliO0df+Tq
qvHhMjK+qo+apcDpS0tvCnapSTH1i/qI+TIlP3HjOnDgm27g3ZtK4muE/7V9jZG0JMD8mq5+8jyD
zUJdk44oqN2hSoi0VfL83Xv5h4h6XBiQoxZ4O5/551dcJN5Zzq3fKZOdC3eRkthJTcZzbPX8dKvu
0IB+f1DV+5gDmzCwIau/9bNMGnv8IrDqu+lscSZfhLyYMdDqcExIiDoV4xFVjSJJRRs0F7RiZS4Q
5H8s0ShTpEFCSfkiYBxu789k9ztd1rhPpqJa55vZhle9R1Bc5FSb6AXtB95OnrhcK5aXSpPsPEO6
vGyiXXGtvrfEYQXX8da6vRRw5bFBtIQsofhTdp9vjS1ofEY3zcJnrfebTyBjJDymdjTYzg3a/syc
3DAD1IEppXulBzmSE9K2CexOfk2h2+WG0wm8LjM5lq1TrD/CC7tsEH4mRz655pXik5QpSz5f4plM
tGwT5Ggj//J6ugmV18YvjkzqNlZcqAjb2YNUkzeZ+Xdz9u0C30wKqMtfUgfs2AMTfccCryJ6AM9o
XGT+o7nf4JMyUFa/V+15Yp8DTTBZorqaAHGndKIgoGzex7eh0kAWMzxE++XWNA5toPwlDyZNNsIF
/Ud6exXCH1V7dVTdQ2a3aPeNxmLj37sC8Cb1LuAFJk9C2rIXRtOCCUVXBV3iEfbWzrlNMgedf8sk
ia4ic+zmnRUBIl+/CUiM2+rGI/8uAv7TF0TIwUxyCjMHhXW3pGw1Job1DPLP+WvOAmpVNjpstuVH
yW3hTsPxnz8tUzTFnmV9vY4kSA3uvRLagzj1bS8g5cqsUvIaLQONGPy4Wn/f6klvsFHzUpOSJcWK
VuRwv+CJjUp7/hsYGJX3mNnsWqO/j5JWpDmI9J5wgM+MWmj4Q6tkyxrkOR0wDk5Nws8yqBhu5/8A
vBwrTtLeD60OB2WS4Lb9W+ZfJP/mL0CmpjOZLac6aLxPIL3Gixvn84Oejaw4+c4cMSCMJ7HezQ9B
DiByI0arbLDfKgb2wDyuonO1ppNZv1Sl9PHabra0D5a9Z+c8zTn5fnJQyoqpb89EXdyJ9jF2Txes
lMNtaUWcX9MtBC7CZK8M0XmL+9DC8vcXG9mnjPgJSLb7lw9zzKisbN1ofVJ1xnOA7uQfCLFCoTBV
bnnOybfobHiuHuGKBSHDrNM6Z7eZlMDUWoz5FbX5QcszizYAnb3uFK085V1jQtx1xbvcwJEdRoEm
MNRQF2RasVPoe91UFqKaBP6RK2tn8f1JzP4XJ/6FYhRuaeFdbi1rBNEEofT/HRAQgs8ba4ufEbOC
JbSk+WNOLrlBnTNX7xiC33NhaWMRSlA2woxBry1FzbUDcg5IDn20niYvD6+efWq+8nwrQYBbQ/pW
G+ROGMWpskJTGq+u2LmlRj+q6SkpvVc2X6tVM+YBXGt+GQa6NK2TETyXPfOcHH84UtE9G7BvtZIy
P02ty+J5gkQ29uL39CoQhc6cXiANUAqDj+tRBVKyOm1KPBzzQIAOqznTk/iwHAXuiimhLyDtcg+n
x/vk7lPPUJQsH2ATDggbEyX6kuUICN5XAIQRWpg1iQjlMj0E/0APhO1ijOZ7ooKNo/MlUd8ZHypj
ONLySaTQc4dfnfnvlscFP/s5v3do1FbMBDrnkHScg1nR7wcYZcYNo7OEOZXILSzN99sGHvLu/6pS
KOiJVbUnZXAARPQjG5yDQvYe9LICzJEZiy8NriOJnXkjgCNJ8536rMaAgTzX29PbQiPfZf1T3Uuz
rwepoYTWNOcTckX+IcoxUaVhOXfyICuIq2E0D4uUGCYUGoi4fsCrymWa+Oo4O73BgjUSjv5UT2Wd
5Ap0qlWOxnVDb38Zd6KGOivjLn+wkVXMOvXIx7f6etz6pFXR7Fzr16tI8egfiYvj9+oLsmNhLlm/
r2pWm06Tsk/U6uGYonwqjCNP7ZhZCNOqUKwqjRkFkQqBqfAlv1Waybe5NRlNxNQ21IGymFdcor86
1nqX3XzT4t4XKffG3d6u8PNS3fpApAVE+WGM/w5efnTPyDh9wRI4qHlp6ZSvWd9pUBYyrDHLZkHu
y3d0SqqrgEyDrokvZRC2ixqoVScVt+dKWrYYOVCnYafP0fBRuZZLNbmKRffW1zVCNtUlerex0eiA
oCVfdwe3DrKVgl1N9EP/W0hlmCk1TMU9xSIrVCwS/T5Jww1/sO2Adj1a9v41xXZwhBDxMklgOMln
IxAgQf0xw0e3T350BZCfHDuD8CsL9dmWw5FfW/KsRdV70MPXpPxdI+hhjVHnqnYE6PSn+Ic7ZJZx
a6UfnjxHGWS4KEo/fu/04y6AHBuEnjYLODMp8QkXETEK/Gzw39WrZC/bNdTF7vLI9m5obyHuepkM
m6nT7a+R1VFwlCnT0/S4UXIdajF3kpW0qckHnH6HJfqNs/ySxU//E/8VYoL77bjKvikxx6l/yaxJ
0pCdILd2nnKqEnAN/7exxOBw1phL9pK7yK+H6LlHPiXTvCOQD5ULIrN4aDJLxSRlAzy6uvDWCVi6
X3XtTOe9/kBlYEkOdwCw7wa7sh5sDYRVjCd9WYtMyeeo5Ls/RElRTx5bPejYzH/4YajOCrSNpksJ
vzP/h38qGOFsub9oEO2VO5cHSei92FH5yDpZvoIKNkBn43msel7NYAjW0UdM2rBRK0pOlBUm0On2
F14d4JaqJw2sZZ4PXPmP9TlxkxDmeNWziwUPS7WOFvuwgMTQTK2WJtxvnnbWDen+zx/i6gr3w+Bk
EWJuCyh99bSxTpoST90xNOTz2ywQFPjYn5oJlfECgVZf7LlMCRXM93QeNYXJggk2OT546LRasCQ8
kSXw0GcSPhMXivhQQZR3c4d6+PGwzBez+YBAjxkyzWv/C4vDYDmO3NaLfVHK9Be6Fqpl9bz1+h74
nsdKUkrf7UCYV19RLNFQZHLyuKko7UVKU8C3TxxnQSYUrt26G92LIQZ9yN/LlR8oqIXRuW00xV1u
sHNKy4O721OUmeaR1GA0kxvxlOpGFYdBOAV3SNGUCMeQDIKuHFnBio1L/tskNQduiMmMaBML/ZtY
A8+uLwhaCiBUAf/KFvgqAVhhpX1SFszWkEhEbQjULgmvR4FW/A7XZrpuboCNIo0kR/8cVOwpoNZ2
Xi63b5F4WFAkhgXlq7EDBeau7ODfHj7RW2279Hp4cF2ujZI5twfy8HKX766i4CBsufZvA0tGM4jW
6KLhXfX50PtXVoPKrtzwiC5CbLuK8A45rdiHHMDsdyxdyHwK0O4fqS1oDzjdzILHPgPzVm72GhTn
5/tyoXkfBABm4k/qO4yR67yKbV/xRirUYG4ZXSQ50wLkqxuLQyJ3cOgmGa9RrYvgHWowBHIeTHJ7
E0E4EsvKjZAf/owgjudphgmaWa4HqPIdRtMB83t8+LMlJIop1lyy1kmci2WpqesBpbK5glz8S3yd
/lscsarsk4BlBnTKymMgz8NIpCZaD1gwOlACtFqF1PguW5NtDBlvmSbur5RVgVPnthXggwNGsjQl
V1EE8byaKf+85AXXNVarTNkXmc/H+Us7Ewd6AQksuENq9u6EIbCzNRCAmyxmKMcYFhkxfCQt9L/o
N4LLlQWYYWsK7BO3+vsHbm/ZIXhNohDEdTmUgYfl+Calqz085wDCnGo1FZ3hOUiF+X1aWzoCYtot
teJuWambYvC3+w0PrK/2WMmor8pl8YtMp8iK+PJ8c5tqThaUQx98qZ+5jfMI9lx1J/51RG6OAMpD
czILj94bTVbYYZ2MGmjbauFnn2GGWUwE5ofPD9oo9Rv+fsdrrvKg/uIMjsuL0MG+6BZaxnT1Xdby
+1DcokmTBs1foQl2+Vqc1PQxQ+KV/cUV6lMPlJDUWFWIQ8N8Dph3uqW9qZBXw5un53oiuxfuekaT
kha8po3AIjwpkNL4GAtahPkeG4HkaBqxl/nW2nYS/OSMA+S+/Tg7a1S479pNge/XZCTZOD4eZlp2
47jytsrOcGZs58ryLy38XpQVnxTCgWfIGB86m7rHDZAJ7nkphQzXrrF7PPSrWJXgdHixZzBVQmjD
OnOgJC9lgmv2W1BahN8kRmi7zaN8/pB38xxVIuddeJku0FhY+0nnePGmYyx5HOnYCmCTVx++sOg0
iIaPwkXnAJdpBKAeaxFW+OXKXCUktoqc0j1W+qf1eP44Lkwa2okodJl+MfzyHZ2vedvMH+ym9omB
LgJ2PcrZMx5U5FpRpn8oGruWq/smOuZpHM10GyQmv/pKourt00hYtiooCKpx8PxueLIeC869/IOd
hzCvukmFOYbSpRAOace127T93pUnCDQ8zqDiw67esFXhw0P+GLEDWwUNAVBhZkU0SndA+ngU4Cnc
yzR4/ZPYpkI8+kD64TxWPCllPZVg8OArUffNuFfM6sJvwbme3QCP8GE5r0YDOgaka7UEu1qhEWhu
rE2920z6CdM0VrvWMmLuI8DMOmqWV7Y5R8EPMx6ovdpdDi/+Sq5Wmrb0cKjmOKG14+KUPx8xABKx
oxX+E2o4mIIGoGDg78dpI61qgyRSiTfRM1rRRKUudmtXCz+v5znHzBw5p4xxSDCdhXsAoWf2Zv16
nixWZCwcbWHA7Zo6+x3ebZb0PDEdwsEkXmSPn5/c6KldD3n83XF99OgwpC20U3H2wj2fvFibarpR
BO+KzAV47Is+cFJ21qOoa+7+1sp8KwuyWAAuzoYeWjl5md3+R9Ok9KpLJO4qnEm9BnJQNet30Vuq
8m2stMzDvjtZvm6MDLKLU65wSgPt5341vLA9mxFDWCJZSki0+2ppCmVjYP7YecA/xEdlUPU2uRzJ
xfpYb/eNdUDmPyx1o759JAogwmlzThUcoG67DI0DaE8ntMAbG1C72rY5myTr0vbOlOqlJq46Sdje
j7fSuyjck2mwyIySdkQvXW3S/oMHVS4FoxUN1O4dG9d9uGRhKMOgdDz8IFCONrs3nKNpG3TOHGwi
VtFqHSvz9qtgIwESjgdIS75lwNbBNNcMNXS0E7IYkxx7Q7qmCwZYitx8uq2PA0X3OM2i9rCSeTjB
IMjYU7W8BwQokmbJouy48zvMm67Ch6hDFyeKD3EVyJw7HBy3i9vlNSuuGYY8F79b7Qm05z4pGjZ6
GZTHXgXww5K1bShUXFaezt+hUddRU0/vnPIipxUopGhYpoBudhOeZQx4wKFjQL8FoqJQTi+ucsiL
l/JGjLGeN+krf1qsuYrEHChFupCBS2/FQ4muXja1c+3yqGN3YG873NNNQlE9d8su4+m7ljxQqf6R
WjXdL5x5iICVpV+AtJLB64JbHmZiR8X7BRNu4Q/kEK2k5WgRm6hOpapmQdwebX90DU0tVKwon9v/
I6hGDTQ0AlDNUwGLHXwuMTvmmHqgI0g9QQ9WZDIvso8j5ha8KxYU4MfajhHrlLt8cJIhpPFUkwzm
NUrQ3qojjPQFOWTumeXY+d1lgKSBLh+gWRH4vT1lHjwYMOBJ+9+5Nv910gPgy8cEkdx++K902Hym
lmfLlYaPwvJ30W8Mr/9BKeA0fBYL4DPIdnUtIYb6Bz/HH4LdiTR+aMdkOMuBnYoE9e8anD6zR03p
uSAPvvA8A1FDr1pBY3upbEevwitBEJnCzS+GhNwZ8+tH8lTerpNKt6C+qiNF483q4l3z/kxKZv6l
ZoWDgVRSsA+rDNcZPws4WNFQBKQoVELUdevPEvfiLBpCMUO0fSXf7+iyEaOxETjiVM3IHmRvxZUR
JwE15isR/PEuw1UGr01P0jZ0iRCQDoMAcro5+xxq0L4XOnLYfS6vh15UxuZQ21tctqtM6Gvw521m
ij+YTSQCkDKt1oDgHIDS9o8doT6/ivY16xT5xJvi/qfEuDi7rbBmCBXjpI2rOSKlYdkffMlG8Bq2
U32NwEGGVTWvEDTUV9WTpzucBx+7bbWmpJbUfKvbGOVpVpJvpn5G0hIMYKpWGlWfL3+0OWCTuIow
RHF2ewikmft+dCFfZqOZO12nP1Job4MqEFd1j7Jp2FolaN1urSsdrCMYfni3T2y7/Xnt/o9oQ0hF
4+b0hEY0VeTcDAFkaFNOA1jKR8zZUQtvXHBmRokrbywN1ZGBK2+a4Gd7G+IcWWQ5GqW+yl1SmDg9
TRxnTVKaL65N5WXbTkjtKIpmRe5DU7ocCU1ZGPysjghB3WfeSBvyXSfZbl1zQE4wAIER926xHTqr
KZe7BbEOr94/MdSJ6tlBSm7I11AbYUyJq/IwAW4aZVEKNS1OWZ+AnSBGXVUjvKSVIG1wgCbLAX8E
C+GWWaPRIwToMxLrLr5KgbFpc2hhNB4pvooz1EwWwE088n5NIBkohWgVA9z47iAb0+ETLwZR2Pru
veSYtKLb1TQ0ccU+VZSJXhdCRR8c9q2WTc5Xxo4cA14H1muj+aOY64ZaiRBmWG1xDyTwDoT6IdfU
JoEgyAOyQkxqW98/Ehj9Eum1kASmKm7NRFKzATww2DUEdmzPC2QcXiZQWucIjuwCIuvr2zFHyyKX
89SwYk5TwIU5iUKPY8uJOlJ++BsrX0x2JPzVHXsECV499ZsgBi8alXJoTV3UhnVC+PLndvPgXcAF
4T41ULqWE7GVZ3eVqslwmaf4LwoMCGyU2dDRhFRpAYjiQVFhHrGeKXyVUpAjvCbV9IvgGGvqOr0F
KAYRsLk7j39TPmypqhzLBmMTs39ZwK46bh+lrIOyqZLskSPVczncczLzk+qDWB6S8NH9lLwk3Dv3
qEOyox8kdsZhfHFVU4WagwBRa1NxesQchu+eGJEuUimSIC+ABBrFs4dRIgxNhk4RGledM2fzKWSZ
gneWhsTT/+aanAZKWdiQA7+5YgwNewH5CRARsJ4hcXfIhHCTPW+Djh9C2AWq7SZnU21Y5TtxU7Bc
fJETMLtuLr8T5mDLWLaogOmvGCcU0GbDRe0fOi61tCe9dyWwo7XcZ23tYVje2f+YMczaAZD2sta5
TG0RHAHa/QMmReFox4W4UgiMGXa3mRf8u/2f6UN5AcvbwcjlQ1ARr8b8O8Psw85HhBcgl8iDHKv1
JiV2H3EvnCCBdTN/WjHryRzsEt70zC42A3+/8LYn8NHt31VvMZAqmhws6HFKry8DMFhv26hS8eoQ
Qj4KAjmqO97/SJtzZIRD4HypLSptp6d5GKQ/yD5hAj4YnOCXK5DzFNwouIRL8ZDdsMaWWHXlEYCg
4j+Hk9Hz/cWNrGWVWaVXgXEHKR5Jwl7KKF5E2l82v2u5SMrpMdXOdLCcMvH68aigGZK2K/c63Nmt
crR0dbickvgZKEYwPCSmS7oOUI2R0ZoFO0IyNnXA8cS9izPK7TQw/UbAbJZA05IZA9jSqT0djSxV
sQMn+Q6D6WnxKEIGPzlsozS5VAatZYIiTaCrwxxeSvvX/hqWrECBhjJkw1TNSLkPT+gOzdTwe3Hc
Xm8b0GXEDrEW8A0kSl68QCx+8m/j+qzW9c29z9Tnvl09ZPW5e9vASoe8Ihi6XItAGlt5XUSQTv6p
9n/Fb6KZXlGRemZkBduPnPAM+1peG6USmYubRni3fauJB9F40eKUiOsO9Ht/oyBiuVv/Fjpfe3QC
x3QGLUjFk/AAruspvkFMmuOiI0I+R+GTgnrOP2rkqA3NMAQ5ULDjBCFqo9LAkhMgTHbeTBXSrLM3
8MdhOVIpvQDT3ivk1njYBdWpphzdSb7STXDpWyXMJrHiCVB966zvoH4BkTZF1SHmslZhm0zZaw2B
9c2DO3MyduT+c9q1Rk0LnLQbpgrVFEsY7IImyn+nXTQz9/btaLhIbXLsT2gY2+RqLI2X2csv9PUc
YHTHeJPkN+7E8m6lulJmOVGwFIm+wVDbODYF24D2W5jXty0tQjo1PusAV1uHIlqxnxz5AoUCTJIR
7Lfj/XxmiHkEzZmHMh4RuIqEDqdq7MWuSz6HBArjfxqyDWWiCBAZf/3D3i2MLzzmXw0Fva515h5l
x46noT0RqCRp74q/sB8babrtxlpe4kZY+D4+0sa/v7CFFm2z+r/r0UMg1htCjsPfSwf4xoo86rHF
njOjvwtas9K2CF8hxTq4/JXcY2D3+XRlqTnEkFv/CxeeN4BmXMUGaFagqLUQnteh636SYGeN2ynY
EH+1nX7Xd3q/VVx8sRm0UjpUgKgbBmzyELpWWGVKPbOONo7n8MF9lbqtDpYwrggQYTPQLSV6TQzX
9O2XLCbHFivh/ieq99m0UNtszZTkXzxz3QaGE22Wvdud93S4q0M22vct3njlSPgH1qywW7AeGBDs
bgBvRh967k33A3SSrPXoFnrSVGd//VjxBf0A+Dkt7A6RcPlm1kAsCJEeyyKdlEhq13oshWNBREF8
nYhuFyZbooIGaQ/BV1TtELOBf3N7w7qF8DrYbJ43n431ecq4FyQpB2DjGbyxqL8a8GEtrKdHorpY
gnQiYSGmcdiz5a6okJVQJx3CWdzJVjBR8ZCM40MtqBD/RJBxDbkpKhhhgs/a4RhJNBY/uJPa1sWW
pfypRVFm+yp5ndNm0ekZ+S6BPkgAi6Awo+GQI/T7FwwALJHLeRXNEY6yUbx3Q1TZhyB0OCpZtTvy
muwFi/yht6KE0iBGrMmtbKOIDjOj47fJxIZqOAN+KM3ihDKFhCvjj39UyUiQCRwiBvphq9iIEo0n
+N36i1Fe9D3TvMiZR4+L3Ijz9nPpufStrzxDAgpHYJR4ynqMK6wtp/kBfg0pOpTVLVBoCNEEoeA8
Mk+AVBbN6aGAUzmA+lc21ASHF/Jvts5k9RMzQDsFRTayZGxgzg661eYCEbeLMyNSftz/O29L6InI
cVjZ0UcQGQ7detpgGEaAPas82CWoketj4Fv5iOWiKyuMyvCP2TtvyRVlxlXD+X/ZSDYaVyGXPwbP
vODsYxX3yxSig78Rc9qz+jYzwEofxdGnx6zgaNXmpAIoX0vElarfZigJ032aJi6wsuMRWpS+szAg
EeP9HYbaDTZCG8MDXUr2EnuM6WN5D2OFB/cHn5N/6yrh9DuDxxffdr3HmhoR5+iUDWdSMJMLcWzI
AVVKeZxPWyMLls/YcHd9woBhRYFS/KGHcsM0i89tweHCtXOSHdpLv6QJff8Buby5ZnvfzKIo+9aX
KzboT4qtiw4wPC46Zcj45Yx1DY1jaKUxoYKuklo29/wudc1yeIX9pUUA+9L2v1t8cHveAvmkpfYz
SIu+mhunaDLgjEyjEsAfIQjlj1sKM3Ygm/RMVkKIm4Vhx5Nu5OV6v5DXSZl85NqL0gbvVl4sNlvs
jCd2bj6RQrsjKTv21MSe6CPIYGHMr8E8bEEl/mHEVbl8W2oyfO0ffmrjxJYSw9L5pWHPgIIgwTG4
TEkAKpTUKXbdKO2xc/JjzYxCXxTyWw77CA48TCxWDYQnxowyT4m2FdBYXTeYRkJSDCtY/2PAvlhz
We0rkzPg35R4TxiToBlIWByyy5rl+yq6cEFBVAslKo9biuhSuwbNjAR6ckZpZgBLt4u8HTi7Wu95
qS9vd6DmCCl251jtVl/MoU/1sFb5bEt97WqiLS9PWFiRgkKuCChAa1Q22E2x7nIjjpEvbnso2W/F
iDS5X5RmTPXrbkdzQKm23B982mwPAvezcekMRJiYJwpdC7/2dIkwm4tRu8MQ5IOmS9c4KDDTv+77
p640xHaPcpN7o4G7/71wUPAMvX1L9WTwTi2vltcn94EmVr1Czi4Ji7Vw5viNXYfyNsMs9SJdpz1B
4VbClDT9R+jmIjIKkkZ7vDiQXdDw7kuAAiKJl/9NzYYTmfaSocBpPLVu5FDZuRYfrWgCFM8aOdts
LZJu+gLfA6yCgF7ounO/uebe2DfXE1llXNOxZkHPpZq7WFRGuhJnoQpASlKq6Q++W4eESAVONGCl
gmK7ARQsb4FtR7c4cCp+59pdfiCOxsdrnfINkPhs9BZzPMm9RAqdd57hKVNYFqtbKpBJOTqJZnr7
OVcaDyWUlANtgOrpaw8BVaHUK3Ojjc1WnbDbxTjkIfd3qbIgsBIP3ocgI+2P3CCc7RpTF/VvLl/R
mBV1FACgsWDFROJXTCafrjVdRih50yabQBgSGNQq89aVpK8FcTm6FPE9o8wgVjxCBVHJH+pSmojv
2cUx7h6bolY4dxs4DZt8hvGxKJl4tg4ZRKCmCmz92UtHLHa4MVmJObBFcs58lvVkyXeHrwzaPgZM
GMxiWvnHmStVY7t5uRP/Ze3CstA70+BIpUO85kZVf5PmKmIqXbYq1YYjt5I0oIzBrZbfBJ59SQq6
2jN6VVDYj5hUHHi926FITWgWgs5A1exde73ZND3pf0ZA25iSAbeAqwYMIou9IxWDu4Lz6B0Wz4Vj
W8RIDDA3PDMzSRChyfGN1qXR8iK0lrgnpX/3rIj03F1fLbNbzW8rwjCCH/RAzSCwpWdRjRGeOS81
HnRHJ9gDOy4PW3bxdYD9sEevDpo5l9F7dRq8Ia24u+8TLkln6S9Yf1vjU7iiVj6lBt4oZBFzJx1D
tB95K8KgWGEQM3z4YBbt9d3/BI+JC45C1lG4PxkCvL8C6VUWXboLi2n03wRgh+uz76cFtEyRBD+9
Czh7TWX9ajX975oPvOFz4zRBMCCvyT6ckZK1HLlo00mw7WZ4KUgMkQyIZ8sPOJ5e5PvYiZQ34prh
MiC74hn1vAcXM8aB2DUHhinicsyMXDp+RvW6VmBBjF8IaTae5CzpisoeZpLzrc6ZuutukMOIUnig
CzYo85QZ9C3alafT2h0bfvWf+Vqy5wwyO7p5fqUydSl1UhB/bLt1cmTE71cGlUfilXoRTdirkOyR
93AuOQNSdQQYbj28sn3i+uub8scdsWCbQIeVoTLoSBo6o2F2kbTVsy1ah0ifNZX6w6wESWZ2o3/F
AE9/CFptcQ/pGDaslCYuztbHzlxA7t6SY/IvaUrAWRcGDQ2Rpkqaad2pBtO6VGmOaGUaIwDU2urI
/K6X39921B8lIyIfgkbWWRJKcBujqpuZVdNf1vENPhspQNLYHwSlVb1btazZ2IZPG9Xs1GgMmUCD
sgIRCQPF47Thbzs68C6CvPI5Jpv/iHtEVktTHzQWUD1a+k0k2u72kKqea+0mL225s/nReXx4kSZc
kd0YfqezrGNqyQD89S2U9Vac35Pkz4OrTOjt7IsPx/htL2H1yxcxTMU00z6Xo/+Vghb6N0uLUU/r
oN339wdsPP+eCMoztwitf63pz+Y1LbTBZ1Mp7+SBo2bn3+PLNCvNTPOk8hnj7WHRFAp9whqXX4Y3
Ect3wZQZ8glYrxjtnDxK/X3eBsGLyEPwd4dan/CicC/hWVrfBpum0tav0ND2v4tBNODeYHQyC8au
nDOb8QMhILhNHPuL+GjFcMdstPhbUJ0VZpMYU14rnqqwjDkHIQtn5w56kFHLnSXPnDxmjgu1Yhk1
ydHfdTm+UFPsH0jW+oij8CYwhyRULfhxM2bhwVp1UQ51DPcx2YBoLGsyLN2xQT9cla2/Arphq5jp
5DeXHGqtUKdACgy5tSWge/BV3/yjNjfQUWdMKMKYjES80Sk62iEVUywQn6TUeIV0XGt1hil+0oJ8
DKoKmh/yrn/ukkcFmUERqh+TRsAqVXn+uK6qw52tuPrqKzmGQ8NTyP8V7JtlDV5CIlpRdFZgWf2O
OiwfGcInHpw92G6FwNBlIrIpEs+vGAMpdkvVOk1Hyy2mgKXFSL9jr9f4OtozkuTgl0xxTvHmjBNg
2RaR+Z4/AjM7qyyFSB2IukKK6C/AGnPAdkJat1N3mHVRxzbpCwBUhucYJLiZITRKztZzZQ43keIZ
2BFAX/bVItC40rsapt5IV7Nv6C/41rkYpGC5LN0i5avcPGXu4My7j3XPE0xghNf74CT6vU5e4D+v
AKhLBTzdw1WD4lbcmPS/6jS0vLsyH6cDhjsURtiTF+xld31Z0M/vTttxdiblV+xIf3R4A+NBl51Y
l0gb37g4ucsvK8y3VM5xoNpZF7N4dIT3LuwiQkz42vesMejGomFe1ZH7NN1/hF4eVlEuEFOKHy2U
D9USk7YHc5Amw8pbMhxdDm9V0lCTucBth5vZPPuX4SoCPx2drwm4CjvIxEORvTYVu4aDgK88J6IG
H4hG2igGovUz0T4oUFJBgxXMZXN7tEQLMqydH6JC4u/NQjSj+KzSD4fmgoBIE4Alt+A/sVMt4ufA
WsTMURU1y7Ph2fSQz+JYykPsDwhVLtD81J+7qdD+fm75b1Dh1NoSHvV8b8PANCSdKEhKlgzoD3YG
VMJ4YnmHMy6DSZKg44yBfqkUwK4HDwT0R0UyLinJfQDdBCEcxSbOeUw3iPmWLc4BVUOJbki8s4D+
zUl7+pfYmEz0DeBmcvICXqLNL/jQe53dbKjNBF7AJK2g0qnIJHU1t85hAltusFZbxrdZxeYAjy5G
c/QoYbVZCstq1M4TAogPt+pS76JbdV3C9aIgvPY1526RjuorcSatDnbvcW5/YJOMD9OayPojhPGU
9s3SI3+03iHO+hu+pRlZNDwFpAYw7KD7t5tSWkhlmV02ZIfMo2y12Ol8AbjBmr+mpoE4xFEUE3ak
8TP5iSjkLEjbCPPuc6OXFJhWCkBeqTU8UTFdHR6W+BFb26784YR0GZIwYrqXmWVouadEZWkwyfgC
7/jmh0uoAu1dRthN85Z3EdmzboDZzz0G6atqiAt40MJqTzWA6X4Oto2RHbt26gf6wBVi21MvRbuS
XE/RGHNBX8lBUSeQ0NNskOJBZBgbP9x5Rbd/3+TuvmDfCs022rgiQFBRrLAGUysOSHLx8Ju1dI2a
8lJ2X4d2j+Y4X2NIv6BqPsvwCX4bufhMYkuEg3VChRt4gylTt7LBUyxNp2gwE8doLZ1BdgpnQkuh
DY0UJ7uN2PhvIJYhZOQffCzpsVtkl943TnwfpNttQwGMl25JLkDyA1lVQqiBpg6/IfVmm7GNxTqO
sgtDxRuwP3CGhOo3esvGhip7hX46gVCqG0X+mknrKDd/BI05sbiWqZ1urAcps80Uvaeh+kUEIDEM
IUz0iSqA2FgBFmz56JE2d8ERl+98yWLpjydjq+AkMx49oxJfDskUCpVaz1lhJvbofTsDUg5mrPJl
n0kwgOSAH+Gut8RamU54g6v3AkVppQ+xoQ2varjN/W3epElc4vR+bLx0tmCfq3E2U2iY8bvq8GCV
yvUBVMjYuBKXq/v+UfMqP6HAIllv7Dgq0Zy6jbqk5vQrSTi6K06zWqLtRZP/OZ8+RrUk8MLG8B2e
lpiAeMtNim/VMlxrqzyXdL0snniy/0a5GFmLKsQOW9G+kjul5QMeNVKlFQ+9QnWq80U34OF4thtP
Yn6SquVLq1eFCrqtp1Ppp0FlJhtn8oykbMrvqanqx9ku7UjPXEzCQYqQKfFmoinmJdKIXYq0WWlv
J/J0F4EI+D1ZatkGascnuJHgtNLDo5xWH9/FR71E6q1dehKxLQAyNzsUNM1NvkyeWgcUxmXO4AWs
+WIB+TQLno5mVA+YXKYk5P5ZUhnp32F5ymObJr5lpRaR79xYzr69Ho1iQDemb/urv6/0edyfN+0s
CcQIRKPftK4aFy2GlSZk2T3Di4mbDlKV/pbAuOFDsJsETNeljqFkVKwE2EITP3S7YIl3GWfBwoe4
scDTCGM8KakCHwn1/8YT/FOn6xwXinZv1lzhayGkfPvo1IMUg25EzlwJ/qQqVaVZ3FkRnr+qh/Pj
FyROVft72SgNBN7dRZ+qxHAHwDublMuKDqU7478kirifStKRbXLe3rFEsN/YrDmjYcPctunsxzTy
zJ/sxtuAHw+uNPBFapsuSREbW5bvtHdO7BaQhXvdKpAPoc5tIbP3f493EZuU2n7T+LFLGOKdfEKo
M4V1V6Q+ISRtIG8DmPUz/dR+RQsvIeFQGBuLltdNAiBoCsTm8Zwy+LLx9WEbkeqirPf1yeJqyiQZ
y/+NQ3t9w7ntnS+GXTDm7qdV38FR+twgzbO18y0FcwjpS/8Bf/Wm991mIJSD/GW4symTC97xu+t5
kHYE6qwHrEvn6P02y7gh8rjNM601trx3vC6bPL5REhRrumGhzNoL04l2m90ZmHPcbbCrLYeu9mOF
qlfCbHNc/9e4ASand5SvAj+OnTYeSXjTNSSJkFKA0UlRsez6TqMdv+Rif5VyuNYr3CxAAftLXwcE
Vc1pLIGYR4F3FOC63yM+/314OWGjJEgcT9373sWG24UrpFZ/zwPAYEQaU6tr//zAyTkcXay2uCEQ
79CTJuZL3JxgRe6s40th0Vz1yQbORvBI0oqSVJ+gL3yKAn59GI6V/r1GQSVcqPHC/tcSfAcSn9Vi
THxQUU2BkEaBw7ue/i+djkOx0463+VlzeoN5Ck0pB4LIvXjzNkN1+yMENuqOoID9043/pXTy+d7w
2TTlKY+8bSypblbjfKREya/BDqrskhbvlJ8jdHzdXVT7153E5vFwQBa8fEIYt1gHN6cm/OQdloIg
0mKvl2QwIFgMvUYiOCC6+Ex2xCCBZu/YU92GbyZaiQd6TmSQqzRaKolDwSvOQ1heGcaMb++soH63
pUboGrqiPHjcswnUchSAfX39sxwUQq6Esee0t4GzT+wo47dqTC6UrzbDdtMxV5t9XzQ2Ey+Hlcv0
jQ14AuGQ+nn01BBvjr9O7d2wsGg+QOGXKwplpNT29FxOH6YlXmfR1v6e9u9cB9qtIJ4u4/CrLhGQ
1xJuYrdhtVdb3g1jU/RpbqDoXD6N/LL0Wvd0J0hjfdV7l1iWnoDJsaytQ6KIg0v0oOJ4wtIBz+ly
YrxCVFFqd/GfiyDNa5W1FTaSmyIGUWfBF9Ig/mnPv1oNTA/FNWsQnwQS9y0X+Vqyg1UuJFIt/ZML
CalNQJ71WZGPLCFWhoaSGGr1yISZMselqy5DLDHSFlEYuC2iO8wBPtumMx+Y8YKM0OKLSrsTZSdC
bkuEKr2wxDJSHhg2LWL/NWFCi+V3PPg9vrXzSbqCqHKxtr9l4sXrviPWjNNdJyLbPpGxotfnv3tn
m5oQmKe5h9pUB1WdtBIWeUE2mhUba2ehG7fCuQUb5ZI5MCvcf9A6R0sVfTrXllCknaz5loIuJ7ZM
ZII3N89uf+Y4XF+tnx3MVLst/8m6JhEYmujaNvKGu0vulE0KPzjoKVbi/p7pqMHWCBzLLKa4XyvL
4X+Aodg15m7HgSAZG9IWrJIgxI0eytcwAUeAXCx/NAsuhmugqxLG3H9OsoYdtCVbw7PXQF9Lza/2
AJafma+pV40iC/9mlKyWb2Q1HGHB35PtZpguofLM69ujtNhMjOEqx6GwL+v2dLmfzvW64mF6fA5d
gxjHuvIgzAmTx0Ptl6jdITcGl4N5FE3uFz4MXjYqhMM5l1WgKrv1s9A0YHoK1jbOWzeX7XmpBIMQ
Sc2+gxNVTs1fTwqC4gZGS488vyjKy+5syArsJ8FJQQmmiBLHonPhiry45vi2mRPOYOMDQb/qCxW9
RG9tbLiqlK4o3kMRR22uq/RrA7MC/jLTpcqszv22jmEjSZS0VPJUIgKAoY7zI+6aYDC8GBZn1sEb
jL71/Xc/1eIKScQXVH4PKCRpeIVac9YfUb0Cjkdqd73zVsU2NJh1F71VWtYM/C9iwN3DpIB1YE8p
CjM/4dzaRKS+8y74hOnhjmpydOmLpROpn2yVW2egpPjXw0rYrC7WpdCNjlzxoY8Sms+MKb0tyXrk
V741zx+PA9Ns7QLihqKfUOWyB6qTyy2UZ2KDZsEjLHjjqLl+w7uHWdJTW2xrKFbSS2igS13JQV+R
g5LUAoBeSvg/9Bp+/JPSh0AyL1YpQUDnOpxHC0RcHWOkgizz/I5sO0ptcRRfSV7uLPurNE4xICmw
zTWPgvFwvv6XMWXPpbkMlS6/wCncfft/0ZIi3b9sr9MdFpFj12NaDEh7wxam3iMqVh9YdqPbcn4M
ovcC1XYC68FJ3ZLnVKCi3bQ2qBpn4WjYHTZ+hLJTw83bGnr4RAjFC2E26AwnKfRVA/MXakXhOzih
OuJt3etrFNKU9Usf4U1O5bbuiOqxLifunjbwmDyDktGz/YTkyx2zOJ7ud4WSZZqIFRwI4xGGiP+4
sWuN3MnNV7bXAYmZw3Teu5dD5JHvMr4XkvT0yUGgpvPt94/Ri7UAubQwAjbsfRNd4ffKjiXYmYnj
RzO+6rrlsoapqT8DpgczAejmdzqzGWTLSRNwJ8Q7MEEsBLqfM9cZ9BYO61nkK0RF1bNPlE9odp9E
tuPj9n1CmENJVIkyL6gQSmlZ0RkFl9VCno3o+Z6LCrQMi3WACmDWPDbfjiQ9W1iMxV8Rx1scRhNx
2VRFvEXOvaRLrt+UUUlzx4DYtDdouZ3ov7MLvmOh8aC7EcrARuk0eHw7iILrnUkcWPAfx3HIzlEr
+AUvxBdfYrs1psoZlfBSdt2YVB/X84/0UExbzyzQhFEYlYIVqmvmyeWf9XZ1/TYD3xQemvXNASNw
6yhMDymcoDcSJPB1JDyIHguSxvILmQx404087hvSYD1mHlDJOYSHXH8i9GPJCNUOjMAAj/8GGlFA
9SZBkfECVZW9qTjUFEvIwV1lqLjjDWMmYIFFHwV79IRMDNJb+pDqCl3Gr7/mfNCxzTRyLDM6qDEX
tUssIqDLprpyvPOqxs3EHFeiUDUK3VkQrjeM3Hhbwb6EOleND/wZcEi4h+IEIIyKNHkDKLofUXAn
mspZEUHdOr3IWkdRPt0CaOsPckffRnHOHg9TeuzlVSEtmCSg37x0IiCqy6YkbHvMmaAAogEFWmrc
Ox46MMYs4aJQIWlHvOOYw1sgILDCbqr+bNzs4xtuAm7rEap/w4os5RyioSwWW5J5LU6eZMGz1eka
T7XXhwLsT5WTdsDQK4cZpNYhw4LavZRkl8xszzYK6uEn68kS+n7Z8fFMIPmtCD//w+Fo4W8EuUAz
YJ8uF55N9Mqiz5TSryVShCKikR9Xe0u5VwmnbXcWF6GioabbEESJQ5EHTbM1hlP1pTrdq+OG4imS
mlj55e+dVVr8TjuibPXa24WPHsNgErv4JmPZ8MImBZhVjmcnWY75YoZkUkZVlQKm51I4rGCqWFcS
CUuOG0JlQpmTyxdxVLNvR/QnGN+D9V4dadiPkF8zhwhDlUwo1udcXlssaF/g6smtdIXi6CIq41LV
/elgMYEwVxz8+NsJcMPkXxwpZ22qV5sJVTKb7vmi+2Xlwr2eNgZ6cul4b8ajf8jaMV02mHJq6Vvk
bAunw0ouBzbwL9AY8MrrwyfvUY9LrrxbdnMBYSDg8xUiHrgd0up1JbGUulBAYMBcvI+H2NRnOXFn
nmVSUv2lglEhMkm168h7S+rOezA2VVeBN5VhNG5ryGaB5EmDIbMYWHjidv3+gQ16N1gG+20VujRb
Hhp8jVRPv0XbCEizZ7lupeDCT58RA+STgp5wOH2/A7GNWdJAbW4Nj1bRRaorVQ9oATQoxSgKLFlK
dyBmC9Kk1lFCd9ZPvb96DkM8XjPpaf2DE/rMFEyY88Osa/ljBejtV1pj2rZmI71QjGeim/f6/94b
MZOPb2wXflqAHu++LXOMOchxCD3OwsYo5KTdJ7VTHqN7UiD45n3doPCUpmSNfVl4gD+/bT//no6k
6HDPIWK/0cmaxXEQjDWu3sqMn3xBRTt+Co2UxYqwU2fhYQfHzabUpoRSt3japM+T2LQhN9QMFWqD
aBgV3/TmY/huen6H3gLOM8TQEHHe0wEN52bFa54Q0dWSFSLpPFgxgccsbXIwPtiGG+rggw/IzkCf
EDGPNasY64ZPv0mZ3jBuS/ZU1BqUwQ3mav+hCPLLDXomW4SmiqrSggCY0Zhbp+mGhcHlkB7anuG3
HM8qkfTrDPMQRJYJyXwseL6mZXRju96LgOALlm/jqrxSoEzSy45adpcyrRd8iq3QLnRw/cWxLX+b
b0ZsirPTHQU+j9VYpdufqV78rWmYpeHtjpXkmPizQfQW/058/SUhfa/Ch8maVIbmYB0OqKWl5KD0
g07ShTzGNPX4riM1DUhk9MydFWqzuwK8Lta4/qnv3UcwkXpMW+oi9SkdtFoxM5/4EgzJxsAr6z77
jIHJyUz9Yd4ys737zgZlMDAZYiFob41t8U5dWFAGwcLy8Tu2Ry223xXttSdoKHjSnswBsPnkqaHt
k/lQ9KqRv2DO1h0qvlGx79EaxzBTszVoy7uOkkg2AJ/5ZSA5VwoWD9D3YFhPVVoShpc2zmR9DT+K
LGBTx/9Dmm3Ranirvd1/GjcLg08dvKH37LtJCrUJpedKccSKE9pH+fD7w3eswGwSMOKoG7OSYJm5
sosyun2xR//nn77N9GUOMmnQYyNzEhTgFmZhY0kuprdQSMHefQUTICx5mKstAt0Dkm2JYcRV+aaD
YAqoh5eA2SrBIjiDD7Xycqtb6JFH8EBsPkc4tHgOwxaLF/IogEloPtXbmMCjdQW2zm45vrG7ZI66
oRpf6uYeLhdA91Lf8rlgE2bReBEp1NoQdsRgJgdIurRBpmS1TDvZDGK7nGDg41kR7JO5Beu4voXG
Ab8fuam+naY7T8PPQ6YYov1QgBmLAvQgkedtd5wSYnfsyBKxfbNPGsnNMA3Z4K3Tq370p2JbWkQO
s0gHRNY9YzgFUAKNOqd9V20JmrZDosJDvGevp0wECBjQnN1qIaEYFhzwJ/cvizAEkk5ILkJ8e55v
heBgiqxRc3NcA2yZWiObPDAsPmv8P2L6k8McqP3WnWRqkNdl57bufKNPX/qEJbd1stYDD6PjpO56
dL9smp1Ym9y24Vud+IJHxz8M2VxkV6U5PZTIdstwGRVkq1r44E1TqP5o6azmmwdZ0Oj2RrnPRCh0
WQCgVjDNI6ndi3sJ6T4tRk98tT0CEiSG2m1dPZtmMYFbzzsUO3VWXaO7J2hJjREAOneq9rz+Rtvu
hj26E7XpXnSj4/WmjBb/H3J3n2VVcXBM/1AAJYv04aD6hE6dj6YAoXrLeC+jHdbxPuRPaXqwrRvr
ijOVSfQkRykdL6aRNGuSlI5L1Xq46DXo2ZoFq7JaozLVEN69c73j0c+oSPSwtulA5VWEvnNlMMde
PR1iACzT6vmNuKweZ/SUBb62N1hqaBf3fDipTKeCfmVghdVKGgLLPpOUBpgsHr3k2lK3R2T7D4jI
XUeQqRAZR2EAbjRrTjjLyLqlzsWIwAlBVoFRAPRLicDCYx3DVpmHoRbE3GN0kTZB7W5cXqZnaFbE
qxixec7XllAxSWjtHyKMoWTinZP5E58Uphd1sDzikdRLNnAaN2W01LjxvAy69I+5EkHXrbIoBLys
+DurK0nn0q3TtXqBFnKjxfjG6Fs4ET1+KCvowEYVSVe3/B+bFMiB/bTCVzJfJ4LY6cQnvIuQcUll
nT0Eq6NEeynj2+iDYQuzk7YLfLrCcYKYlq3B/9UeGSsp0+SBNQrfe2DsBRZfFj8elx0CYS43vlge
1xlPvwlVyqJzLWwVqHA+vNFaelg5U5M+X1vybh7ENLwWqZ+Ym2zLj+25ndpP5DUOIlwMZZr38REW
N77YbGNWzjF3gHN0tarRe9w/ja+uzjDbdc1YzcCCpDWf0WVJR6DjvhbpzZ2jYqM07iAyI8X/KLOX
IK/dtgGOAo/JNsq19vF85PZioMGSAWFONVifPmoU15Quixd0ejNxURXulBMy+JbPh20tpSTcNx2z
/ovfbdIS+txg1RX0BFp5oQNG02eSSermATlcBnBy+pVGNKAAz9bGuftNDA+tFWzkYw/zfXXY4YLT
9+1/+Y7J0itDAd4zFeJqCTWisojFavNjSW8xChFkM+YMVBmrr7jHJj02CuE934cJfqpiUxh6FC6z
NLT16zHxHTmePduC7zLMz4Lsk63iN2Menzx/dguYlJnYs5ttxT8vIlzwZlwMA00SFuXTjOKYi4ZI
u8jTY38dguWdEYD9i71kMcP8UKb5YuvDFPyW3570roN2Dd8EosxnEj85WJY/bpVBW/qtpLh9wQRG
EDX0zsy5IbrmAxEnUI+KsXZM7VuWq3YgbcCcfdvuL3lmcV8aLb8132Q1Ige9K7SnHvA/WfPBtxMX
cjIMz4mdnZIXIOd14VTGcc8skIjW66KpAM4I/N5lRYMmBBxjtnNUkaM72oVMlKsJAdUEQKBtpbJg
eR6DM1sZ1YjSNAgeJuCLcYk3u/pfQZkaZFqfZ8Z+hSCOoMQ5dr6AVlolUKT4xOt5pAzcPPAxzX4y
4TTd0qNGitu5HRs8lIN0IiNzNRE6i78fO+02Mmll+tSKwvWujQlC08q0T+v/PplWkdZpsWi2HoJo
CSEHRSnwwv5I/DRp3or2hIzkaMJ8gSQq8qOsxWLRV5gQGRbL7rW/c98VTdcOHeVLwha+2RhPMsZG
h1TPpSOFakR2uSn3I7tFnpavjYJHWWUbUMt7Msz60c04ZF9v/gry/5m7GIxqm0Iu3totz0bvTZPn
RE3juPy4JiIp9Q+I3oNRh6lhdrxHaaaP7Xh+4rN822/3S0Q9mW3mXyKP+JRrWZOvA5MHzqVXARPL
i8z3M1O/Wv1yIWeCvmsI7zM9TxLPgs1QwuIqXnsSu2kyxsKXl83hNSq0g3CLALQ8hbpPMgD24qK3
cHf/TEzhJlzsBteKQ2sPa9QpcnsAuPNx51aHk3hPqCRG5RskiSiqVpASFME6a66l+n/Os0I2/84d
ft3bdMG8YviFti13MYj3PFicN6s8W1UnT1qnNtZMhjtZE4vuKoyhpCqthCOZhAg0VHW2gtNILGft
soZfEyMPu5433q5M+ZQ3G33iAarJvVEfbVil3dCUqtkeBkq2B4fzdWuLGSnLDkigrxIoGmFB2XXI
b/qPuCi/YepWhdifw5x/IRTb2028VLnvmzxDHPbfRuGl1hoGeQU4XdMU/nQ3vt+3tf/xuKpLWp5Q
ZI3CJWMO3fySHlXVCEOqjfPuHdTXwCMOdlcM9QdHj5aIkIUHZGXCRRFp3/+GaN6xQIyZVmwAkQPr
/9nS6ILf8JRDsD9Ocec8/pF0hStaLD+4Ax7a0TPNpahDjO8Fim/oEqcbT6qAyLf/sEGH52N8/y86
vhwwOLUMU5W/VwKoL434KsyJNmmJFGUgAovayl+c5A3BSIhFWBeKtpDR0MQHEkTH5Pqz/dqbAK1K
VsJJsHR6ZrspV58v/mew7rUhFI7Ql39iRr6rvFyYfeLW7cCm4OnF6MKfTTcBqfdTtJPAxml+eRxA
oOxeRQcWo2FgEOzhYMGsAq52oOeT7AoObmpHfqWQawbFEqaP+j0FnMC3TsRpWrjlB+P9YymAYYNC
6Hz032JBjKNN2xjdV1oTlHuVcFsdSYboj4ZlZ3p8UtPqrYntGNwjjCF/SslyZYSX7LPE2DOLw332
EIsPvsMpKuJTppZ5sAeX/mUx2OKDh0no3Vo/AT0PW3WCDoxLW4DUf74iqsp+X0m+n+5L8lt01drN
Wb3BFb4Q14FaBSDpnVP38tsXJptmdU8fNl7lOcVuIOZGhkwxwmPi3+s56GeQgrnrdVKQqTQ8s0E5
5oiqQVJZn7AbLMxvNPc5xrDWE7LUfNaPCJdonfTLA3au0+DijUtqbm2AGP9qZuQp+8grhHvgh5B6
C6+Rl5YVtNVoygT2F5b6htxl+C+L5PmNmFnsss3qwgCsbIz0Cvn6tMnvHoUb6rruTdHipnSRU8hu
5mHiwpM5pTTojuNY/MCyljYrCIouiJO9yjqZgLKauJtH6RCcCtayVy4Htb1v3o/EiEVLzmh2YytU
JVeMoD/nS9a/Ez/zasXW5SJ3TWDC8DFQgsX/asIgquRkDebnUHc5kqCgzUlIgKOtJGIxjmb8Pa9o
U5p9LwZYjcTMXaSANxUfBWTZFRVIzL2OWkaihW4iqGdF+pHzB1paVKb4sJyJ3SYtOp0FnENBsggh
OeLBwmUN8zkB0afOOeNffkeXFklEUpg1cyQwrOCE0OQ9whEL0yNRtnkW/NEgRzoNesEYuQ/Mgbx3
bmZShRG7MqyZylWVuUTKUlDIUzm14pGbmTp9E5f4Mdkyaqjt4qSDCa90vuQReFHH7UGIO6hJyQ4E
eF5Dw+e7P6gdmw1XaFDGnOWNcTEJ8fIJ7p6DnJSbn8fTWDK+fJBhC5+KLhY5inXWO3qtcXHmEh7h
Ad/U67Zm5woxFPTguJFc+3P8qXMoSgyQTd86yY6/7vs9i1Hx9M2EvqPkNnQHbw8e3SVGEV7H4CCo
gWeY7vX0zTcbaRVzazdImnSQC7SM9ul0zZZmaw9BnROMPNgkBzKepvyMwmvYjdrvkWdV/Er/2/oi
YSBcDwS0PVx3K8AUzaWlGd/TxXBpDOPv/SOGmj1BNqa/h7vB5p2HSeUExMkM6CKlKnSXRx9mJ3yo
C2N6YPEz3ayOkgzAq/W0antZUu6VCjylBkBm0oe6lRcaGrYAbi30QGbLtcTUG4KFRGvCNan89TI5
nPpPDE30WHWFahx0btwzAAlD8ca36bRvb2FbdcrI9sns8LNqkTl591nMhEUkcn9QrA5kr5810qoY
SCQ02HFXvQxEXCBcQ03r99+4AQZJufw8j+s0MNwust+RvwXnFRouTlp45oSiUQBeXvsSBzyRL9TN
R6c+M2KIhGyTCtUFZcTVvkZEMwaXcejDPK/ewa+qYkjBOLSxqRJKMRkOR8+opsv+pHe9LPTj+2l+
H3meOntK7+8cJRW3RaTyqGZ0eqAmItk+8FE9n0aOotHMY1wPQ9sJR56vnKRsugRFgc5Cs7ikxDGW
AnzNZtu3z63Ft8psgTMJMTDmBhdfz91psDjaUlJqOobbvAg1iqJrwsZcPy8EK5lqWbINlJ6y2i42
FKE5LZwz+Znui8CiFcj24astepn9mXtDbuAQKlcTu93TZvhyfht0YJ56goRuOmsoFdJkmWfHW0bM
XzDOCG7O5rhnEEuJjuBfxaCHrJOujyQOlUbBpzvZsFLz98x1yuyxzLrov9rAuyktRlF0CdHLGcEr
1eVXAGwHUISYi0iK7sLDNvMEgMOK9mwjB8a68B/F7+RJ0HxA1E5Lc/TbxJ9E2x1LYqSOzsiYsILK
A99D+cf6MHdv0rbAbEQHMLbvUQG2zVzPboyMeO8qQQvVMAuklG5Yk71vGwSvdqeakmIVhMDscqFx
52+Sc6dHqdOVDBaekOmt+5MW6LcGdafArjiSuC8b3sHdhOq7h90VE94kPgS51Ro9mzgOjkHF2ioW
T/KFhoUsaJ1X1V7wjpMV+nqKPKDvCshfQTQo+HUcRunQpYFoRz9yxe4Y3CBFij9oRtB4URSVziIz
+x6mYjgMkJffmCH0M7xzgfhoaIhUvvqLv0RPRzFnlxzLwb7Nbp4dbH240HbAs4rRngb68TWMzDfe
v+gTVTyepiwRp63lzPDF2vSQxyG8NuEXqUvQceHHNWMVWKVcPeSAOVE9QGt8I9V3TiKrRcb2cKqR
wctu/qc8oMOu2hJ/rZiNB4XEdxY9uOR6oGKgE65KIuSxcV2K2cungoVtY9WjAx5VVVjDt5YhFr03
WxnNOSb2EoUSgXgIhCiZ316Tr2WSRtfCTgt8Q3KUgV9+RlM6X6gGJ5aNgngXoIQK7Wo1CcGBQV8Q
fdOPui691NknUP8e8raNAhn6vjBf+jajvgifkAbJT2KHIlwVD70Dk7TWNdDs8wQkA5gfXC8wdQHh
NMDwmXdb+oO72I7Jpa0ew3cfEuZSawEyKX8vqeLb9L2MkROzx3Dk54P8OQS8wTta69IAIf5C5t8E
/Zun+fIqUmfZzNUc+KT4+ZA8zkkqOdT/Mkf4PLxjA2pF6pRXbepQrrSyVdF0yD1igbdMbzwzXpll
UxMNsB7ig2z34KUzCJKHZvc6fanMPpc/e3HBSnj9guysjeXUS2ve3bmPXYkUb78Jm/FXtAypIihh
77yGm+sKdbqbTb+DNfeWGuYD6JbwQs7g1qNkGMiddzUU7o6a0Yf8qyMjtR7PaKn6AFFpc9nVySfA
W2ILPLqDvYX7zsIadVmUby1CyZIgJosxyCq31aaitdhloYpkoMOJgvv1tc39f/5zBUhCUBwOpTdY
9SD/MB4deoU0TuNdPj05I2VAaKkjGMsaOF/hC7iK3HQc/2+oS2lP6gf6SuA6FpSEJmXTbLMkpU4D
ugGbJYr88YGriv0m6GHr2yLtyoUw8Bk3AW/k+zK6pu62Uo6tAOQeDUCoUThP+Mk21OKdzmfCSc8G
+KrQ/XZ3uugwYBMqzbuLfsREo5COYUHylFdMxtqZGN+3fDX3lWFdU3sX4yQRZKFIh4435iuDfhWm
LARSPX/HYbIKQwR4CTkiw+UBTnWMbPMJkB5Pj1X+uQ2NEbc1ogxsp1kCpqn6JFBwq4Pg8Eo8zs0h
QcarCYwCsXhM5IbpaIIMV6PQkG1bR4cMd+KWN8uD2PlABUkthbgbJ7hqQOvR3kU4FV0Vs9iMMi1q
/zrnirB9xtqMb+HS1M1dFAkNw5jV7Tbxsr2ERxVjywNnmyMRkwNK0CVywIcqJaQouHhy0PqCLbVK
gyFCLr+E3k/t+P8j7WL+aeR3r5rwcWx91zKPPf5D4aaPZHpcGyB/GrXdOGoO613eDfIUdgFqFoCh
czX7CXU5wysmOp6CU8lNWEI51lhD9G4Ax2J6Tp8ly9v00nBpoaiUTbCgHJZu5n44N29+sSuO3Bc0
v2e3rr4fOl2BRSk54KU/LisrpmxMkmiS2ysEsX2Nt3ZPdvH4i6aQWAkLw+6nCzGCWUOtdIdjj9im
+y/vyfzweGc9sWT7+6un3RZOAEXStHV7QWjLCSsozQDcmYgA93lCEVG6j1CGgnbYvjP0NF8svYtZ
N26zCjFp9pOD4XzTXnSKkp5oxB5Ah5DNyRCeHFPbssYiVk1IuuRTa+SetTd6i8AlSPmkDIr5OJ7w
C5Wc11rttft5cI5JyZehvUIvRUkZ3WgQ88zqvA6fCTuxelqX5qgaBl6Rg4GRa/BaaGyHk7TkqPhK
b+20z+eBHaiM00pIIXtVdzfgFoOjU44+V41kU00PauYyvF/CIPthCjEMeUYvjF3dvtMYoFb99+x4
7KNvD7zN9ic3GIcpZWljV86044dDaxJitU03TwLnAbp4Z9DzGa1JqqJESuC+n28JBpILkJX2nKXb
lUFAl+ePUPvs+4GfqDNk7ea7zTozeaIXKcQsWAuolM66124GIuRDLwe9/3WL36L+caLf8qtef1qz
16yHNTxvQ5PVUYnlQt4lT21FdjQSNuEv3KIOQJG1P3HVxfgirDA+lSoe7VSj+Kua5MM+2ab4ThyO
GBdixzxB5e5LemggI0qfeCewlPvowx6ClOUf5tzS2AJy/w2IUbC7c7115FlrFiMUnXbtKQGQGejs
05fzHk4ynw9xlpce/hfbhFeCdnx29oo7lcEhBRpzNhz2SvKOVgmxCG8yvD/FgS9cWCJgZs2MWrtj
+0Qi12FWylAz2IJ+jxqNhsstiAcj8KOeZh8cqjfrnCNUijsLTqEvWj/D9YmkTy/cYKJO+rdEy+CE
j90t1sfyV4yhzdJhYFwDv+GjjL/g+C94wkwTQX09i+Y+8/yO7EZDvWluhCLGbWuzqDyDPMFp9n1U
U05PhK5KzCuvjQ4hBaR+VGhjSmWC/wk4Bga0hBB5GYFTEL3GHE8AnviLDiMrvUmGaoFUCjnoglCJ
SzdLkm/iAQCdjhHVxG6CiE2DZDEpE+i/2/3bR2CBv7hiyqNbC+MKg5pLSZh4ltU8oAiF/8wMJlg9
EPHAaqA0TLcOBJ2mxhCb1NMZg28Y2i//qOLfhgppj4bkY0y5XFG36h4ch5YAo3/BElMnxCUoVFqk
RO6vK0aX0Xmm7ghBfIUMyEIt4o13AEUSdPeRuqaTZ++KWpqTEnm+/jsBCkX43awjnZAtO+htddKd
fezRxWinsLyOLYVwR1YXMqdn6dMIBxQ8sTOxvZwc0ZyJ6N/qhAqIL984uouY2VamkyYSc/ulPZtx
ZJKXZxsk2NZ/vEUV2ANmE4aTFKWbkspsgWKtA1YGqXoJXE7J/26EnTCb2jeLZ78JRoSG5Fh1zhKY
efPpjXsIsWl0/HX6PwlKPHvpOi6J6PsisN9A6rlUnmXzIU53rQUFIDNwYiZfrzkh6mlvizXOHgQv
aAcN66QyGWrXCaTU5yUGGAV/C3HNdsclS/ohakvsGFwLZ+BXBjsFquWuYrfc6rgTN7eQVW0eWWWE
+pf4qwyR+NbrWOijbvcI8wJeIcb/pojLx9AlD9pm0JCK1Y6z/xKFf5x0stQwMGQPIO0ny6v29CUb
MeRpduygMN7mfw7fUkeF4+M3XBXY0lsipR+xqUUQjwX1ZXTusoO6tkKwBwP3KWZq7LcYymANVSI7
dWMjzNmzKYUbdUVA9j/AMI4bTSKABi4K0Hf4MQR4LoF2/pBmy2BlSCNE7qRO2QtcYAigmeADfuv4
SbQCRP+ByBWs1i/8a55eiabjs348cO7A39HWfPO0xbUSR1XYWlSvaoBkSZ0LxXOIEEmpgnTJFAFR
czr4Accxtxly9nKgK4TpVQWYZ//mmfNmmmvH9jxH/xV8LSfpeed8dsupw3N6NEeqp6QPxc58Gl1x
UId0BsqRVb+1qMPkYjK3sH5QE7GWSr8GAAn1de0QldkwRRzGfc5gEOa4YMN4TN80GeLNaKAU+31m
Zfj7frhXmiCNlovvk4zY7trPq8UQuT+s/3+rnxSakXVaZzObD/Yqzs4yVkUitPd7oBhnp6HcvhSh
5rrsC9/g5StZWAJNm9HEsMgvOA5J5lIx6f/q33HHgdxXNQA9aOqh2x3pFJ2BhA4gaQY31jrtcnDa
BbjADTB3owbDLrjJyODUmN/I5+V4kTmACNjKk2oZ5evxqiz6uJzdiu6K/bnPQVGJ2yXXhRkCePjj
JvawaZfBLwJ+No57LVw3gR7lZ2jEExyVHM1nyJOVWiK1mwLRh0kTGuZfo0M2IdZzvkoIU5/exMLH
lbg6i8/Kvy+/ObV/i8AEO+YbNO8M59fmsT7bn4CdQ7QwXcPSdjFM4qiX9SpSH5Rvegg7NOcsmWR/
7fgnPuoH/4ZERrkzi9ODdl+mkngu3yxnPhWi12/CizbNNT2jnjQz3mK572FqWUrgPfKBgxwfpcZU
vp8m0FRtMNrjRd2d0uSvaRXrsD832Dth6vTFRDvuvToj9EBEiE5G9+spjawAsYA5lJxcjjqno63i
TSRvemjldkoILkpQGcJwOoH255zW6KDdoDJp2wWk72OxDWKoPqOFsY8Jrb3jLgSnTeU+daWBp/aN
UofosFA80EtBGqmP3wQSD5c/aJqnf1k3PcH/riDczoP88rxWByKmquRjONMOGMvDmES6swU8993z
yHr+twIV52eU5rNe5g0e0lJO1uq/pMp8ErX5pJjPORcuwgXSHfzBYrcWCl975Hpr+aJiIpVjWuuV
pN7q71xW4Kjf8eZKAkf8ozGyb1t/jBPjpyeTz0kjjwCLQGKNuFCv63kt5eiwmqryQMCxPsSH8x66
rlivBswT4fpgLjJPK/MXg/R+P4H1Bu7ZZwAoJSqltBYK0fMU15AukhYZHEVUY38eoYUCukyClgzn
LW3VO6rYTBCYqNyVvQImFeq2kOMkxk7CGVRGQbfG27h2a5PfrMsBzn1lroUCDjHk8iI4ZKhOELCJ
goHQjvM4o843DyZCXrh5LkcQUFYdGAHQp3l6XG0LHdDSLJPBgRtnMQBuh9N6jVWDbFoJ6Itz4SSc
IQar+W1IAmepRx2Byzq46s8FRvF6UK8brPbNWloQABPpVGcfS+HlBqd4Lgquf9wn5+b9Ih8d56qb
ngE09GhMoZBMgEqhnAjDozvvPn12nuoTJxYU+yb5w+yz5tnjT4w77IXoOUXMVs5tsEqZNb2kowYX
tFio7YRWQ8LMnTa2MQ+wKOUp+eXcwsaqaPgBnjSyRqdEz/FcVXJz/LL+3Zb4YpNVSVeuCkC2e2Nb
oL8gUw9KlXV718ltQbR5ZG9oglhxDadu/KqYUehEUAfWS0t6kP1LkhTraxPQDMHKpPBwg/PLUFaT
AlaWqSG3B0SUfQZd/6Hz6UDy7Ags20dlNM/1mzD8lzbdYl6yt5JonU75IddM3YLl0a4SQ8bYl1u4
t5KcdIvnuAb6FkUJ71sBjUT6zGbO74ce62QzahwfweHzY4XdNpHEqZGp5CHdmoqF6aVofo7KDnjM
ZTLgRsBOac8+jSYGXywK64ealZybvotFyHwdfqUPclxiYYjQZU97CjkaV9EHY6IDmYzBIksosKDX
UPSkyObH2uNWEmf24wbhTr0yFCDDxWtDA0P8PLZddqzoYs7TkV4LDCrOXFBrF9eK0j0DyVLUsPY+
fhXEwZM+hVmxyFECnQAlGRuqIW8F2TRgCoMUCTpNaglztnCuxh3k/UBXazKqC8f8kahsJbabX+s3
iGLeXmZbh7mcnooOg3EWUBaeXBUGBjHjx6bGCjtXpg8P8mhbXZ9Eo/oyzMoq8YQV2qkOPLi1rkFh
rq9/Fk1nl7stV5hONU1eS5YxZ1m2jKY7rPe0cCoWvooQ0lcYtJQigZP5L/Mq6XZiRkH3VEuS9g2q
H8QTUR6BZNC9S5ENKtSqMa8eGd9woinXJAXwKhWsDJs45kH/1MOFR9nFl67KmcmUhDjeMup5ONNG
HpgKjzsrtdHQ86Yx/UsQBQ3SKPwzPnkx5MAFGF3P/m6yfUyhOKDTrrmbxruCFdZB0Mim+lSdA/ix
PXs9P7kPNle0TUQZh4ry8Su2p3s3sLCfHZSO2aBUeSbd+7tZtAV2OmPWoPdt10faC2OJBgTP3x1w
NOWb8YCkepR0fSnri1xGTd7eZwtOI3lytO4V6XCKV1tjUPYK9pRiGOLyd4lGxjKVEwS1kYeG5Upm
z5XdFk23omdjRGsDiWPI8XIsfa4E4U66uTS9I4ruGNtg2mYTpiNHPX11LzrJeM0kkf2bb6Kg67SV
/K3Hz1C0KW9Lf9lfW8fRLMMc4EQoJTasf2pW0wUYEgAf31F6Spr2J8ja5stjy1ETS6g3q9jS3Mr9
Ourf/G+99obUlVplQvUTfCB8VQaER/R5CGtKuZClLT9iY7eYAubtoKj2ymPWWokJTlGH1ft2chmA
605QsEev0NiW1PqGRmdklD1Z/B2sVdoy8G0B6B92Yj35UbO3QgYVHpZ5/CQniVQrt4CxNyB70Qjz
h4ZR28Sv7J4+OR1sl1t/p3rLCxJwabG4wRuG/LqAQja8sNoVTBQ4cEPI5GnE3PBN6l8Q1xd6Fi+p
JUo7X2ywzHcjuKW9WBCf+kskNmN9SZDdVWKfSDCnPQd0V7X4H/2ivBC5t3HM53iLqS8W4fg/W3AO
EuFoQtN7Bz6+3llvGaqyP8W9n+Z0C5LQjv6tgRmE8xyAwe0+4Su5Y5jneWuMk2z7IEumV/Vkj5IN
t+BHkcDWs0X28t1bb7VZArZa5F1EBcHjOikfH5XPaAF0EjiEJuvPxDrw/tlLYesQQ7uroBwZFvnQ
LW6+vrIMHaeSiA8DB9iilzZJK0dH7tRY48QC6pstGSfO1KW0Dcm69CngkCrd5O+u1A4bKI2k51Yy
44sqFJDWi0kTK8koow+FjSZXK9LZ6MYH0yU6IJ03llE7Ww8FtmAIOXMQa7LUCiqzqseVmwklQUH4
uz2UuLyjL6MCcYKcghNIMt/w2WK9W8ayghSR+B9vOCvX1PWApMWGOWBSupzucgKfOVYbf6hi6ul3
C8aBLOZc0KF4Lk5wkF4G46oEEVae5NvHAKWtBNOZvzWLYV+c8lX9KefJ9BpiZoEToz5LHzyhbphU
DGTi0P2fAQwj9NNjipm7WWJo4kzKT51JB5ocsOsimodolpgDIu0T/+jOxftYrC0ERdSHD0FIXdjL
0tRm2HRXHDFsrhBjT+PXjDVylUt91VU2nZQoyzbp96cGoiC0KPAydeubaJ22nAOHxb+huaygqa0c
NuB/z0l3iP3ysjOaoBASY/N25/Gi6FhNvkhmKLQHnEv70VGQrTsM7Ee2beVqviYGulpvspJ4QBzD
LdLFS2cbTfqxOe3xPLzbMf4avr8xx30tmw+iidhPsca6JdpvXrmUDGkFLonLVXPsV2v1sNCPm7+s
zdzicOs0fsq7AgK+CZvS5D/ibcoJk/2ZK3D+17eCVMIgbbL3s434kJE+CB5FxQolFp0CJs7DgtUL
EHaAYCYUEjQUFI514WgFgsqnAvTFYX38aMfeqUDdcqEig6orugyeg1pA/zYkOGVhqDXmUJSQoUM/
txFdz8ZG956TpUJdbk6DCSZf9gMSxT1H9ZQmsCQIlILHqOcY97XYGQPFmxKNHlEbyTwsuZY6taEM
5IhT3BHEX6DUVo/Dsfzc4KNDtdQ5XQPXzVbotruKK/7gg84i3CYBEm0mIIquAJPrJ0ZwWtMezM+X
aQHOALUh7AhMz52aIvvAv3kVFJ7Tc2G6/5b5ZoAYCtQVu0a3bUndKPiji6o0eHwcMxFdGOZJ5hq4
32gihCmYRd1cGNbykEbsn6YDZRLTAWB4vEhHcBjAguGvlpSN9W+/SxF+diT3pHCFAfAz6CZ8epw3
w2w4W9qDA2mINL8oWoIAI4xJHFdRsU8Mk53HgV8RbDQgodL+5hX1L6Tale5tywGmIRmrzI5uSyOx
9HxKYO0K5QzSqkLBPAHg1Ae3/5Ul/YCA/NzZm2xPtc6l2rwVhsFMkNG1nyaSh+hAp/HdAe9qDdoU
t78SY6N+ZBVyJHTG/fSms1w5QbbGzpFREFYslMYhy335lZnzbs0kAVrKfQ5iCW59+EPAvaQ+RNkY
vWw9bq56S6xTwp1W3mEL5rMRDZGzTen+ZdAtMr+QCW5EAzJ0BiSxKi5dQzrJgBAUe2Pa7fRMkjKY
T3efBpaqNSiDOSS4HddWhlG6Xgzjsm7JOL1c99Z556UYMMUe7Lh0Tujev8grD2WeWfKc0ZoLCtoD
YlgmrC5wo39GjvdBluInJwygAeldtj823bSuMfbRsOyg+w6ESrWfuhTGdjkIuh+ddW+FMhTOPrlT
oxJl9v9dgV2bN3QSEf+rIZ/BrecBppK2g1SvSo/blQxqRxO/QAumqJE8asBp/m3gTFjfakMV63Eg
YicR3+q7VE/pbW0IqNMz+OWUN551N3MYqr+U2bUOvp4jP69WAmMfuADO6/qixgQl25gmBrH8jBvv
iFOpaWTSBBwCMlDpiDigxPMPMTM8FO0BquDiY31PaqXvz6sveBJnWwaN9q32D8VW+n2Tu3MHRmLI
q99BpKklVs1P3fSokrZrz8Lm2gqrZBlIonh5yYnTy994ehRtPkbg4oG7rj9W81QgyWCcQd+2LB6q
DLi3JmeZu5s52LsRBPpwJvw6Qipvz651046tWPkRbSRQq6iXsvvuZuXCyMGf4yVQBBJlNLJ5mFhI
EGkUcco89J7QSi103kk1VAbkKW6u0OUVfk6m173q9qM2hJH5KnKq2TcrnvcVZ7ZAlVMg9yxUeKWG
II+50HKrxxhxdmEoUm2Qc4RFZNbkLci58fd2J6dETzcfr9FkXZuQsag4hwh7CwJCzL8QR72f2Y6C
oLkUGJxudD2JWXM2AVnvaGd/DfHvF86N2HYuQIwNQxlNjZ/ZW9pdV2SVN7IDg9SwQOBNMtVDAgCQ
BZmp/5og1NMxvlZyETTYHwBpmqbyZBDctrFug/Lso/n0uwo0uwKgVn+WqPKlm/Ud2ML3zPH7Drbq
w3KRW1AQ0Ob8XqHv0yJv7+2mNEeDprWjw+T/apUXbscVO2ckwcLcgNMUe6gUiwnW67HEbrvMe2rR
4AncuUP2TKeeNAtV3TAeGo3vIPVT14W1GzATWcVx5A282GpQcfcusvikCr5nECxwY8rR1kddPJcG
ViKObxX/6nWnvyGEfaQv8zv5hYG61RWyPfVpSAD5GeAsbqohatHeZbWwQ638VuBgAnTuiHuh+jLR
vUgSOrCq+uyE8hjvFHgDMeaV3gK3CD/7mMoKEBQi6Hql0T7QocVmrWNtrfsa0qUVRabKao5x5aQt
prnKzc3LLSUccEigMEIN8Xzma5t3eYgvitDF/krDgEoifu0CmxO7+ivdg+NOEeHyoNsWTy2H8NO1
aHLZZt7jgw33KisZVnlw4PKybF5Y+zOP7JEug/TTHyi6Wi8MhPyp8+A7KJLh2VvuXd6HW0Wo5ur9
Lgz2dFJANOl91fAWBuqTuZOWG19B+mvh5aphydBXaYBm4uHNPQvJBofL++XdFzYbJN5DZ6mf3TtH
1xp0iKQ64etnjah539hpau/uVsGlMVV7kbUg4Z6afEt8QpBxIh4I1XcFzC9z4kiVeFvWiBBJ+woe
uJd+D8J9OXladHDLTtbtfAcyd3xo7cHxf6GO06qYw4rs7MsFQBeVrSDEUkXbIYgvLWTmMuyUYtoq
Dm3A51TCbDPMXd/j2V3R4k3zQifnYUUsX2JLFfkm2wIfK3TloHR7mvphNxZ0uAYNaq26aS/u96fp
wMnrVb9yfNAW/ZNb030xwF0vFU1OheQvb2bdN8T+ERvA+DCTIWTssRmR6ha0Tl/fITCnpBCMmx7t
USPpm0TT7YgD7kwbYqbxcCdfNKtx+5j2NhEESqvo2cOKwenKbH6nX+2YbTuAbJxOqNWMPH0V+8oP
h8Hft0vy3qwQQtiD/t7oMq14FCEBS4c9dPl5vCPGlex9UjKoOO8Y1GmxzJvI+oxBLCJTuthJFWsw
fGQBUEXb5NcD0ZJoXoelwKuds6kpR1SUUtKeOvhOXfyYHLlNXj+Gv8Cass27Iw05XTiJ24mKW356
DVeY8XBiz4XGxYKPKF289HxCDtImT32MmPl2Dqpji8j3tBHf0AAVVivi+8Xb0H09WSsF4O62HJEJ
oc2Wxs3NnlquLin/b1QgFDR2dGL0KvzpqqDHS+chXF67SCu19sp+SqdqElhYS4BYiqUWH8hGAktB
JPfBPKjEfGWf8QttUsWdEK9L+NEfnX/Rdmlf4NpiPvMwAI39mh/9BxvSdsnAvhG0OEoovyNfG4rK
cRahtOrEGvis9Ye0GY95Xjv7WRWf4uaZIZGos9FXmxfK9ePlETFR/Qby/p5XomMochwGzTnp72/p
DWKXPHC936NrfDcltR6E9hHVCFdl+xQaSx06PF5fmHGCqTP6zerP2Jven9HkSyrTQgEQuq3BXkjG
IW66cdy+N7QXKzCqtploLlsTCHaDAPUY5CEalLxCDc9hsxZoayqDZ8RbCAPLFEx0GBi+MEbiLwwA
FGLIOEgDLrTTuHWARZPcHc1gycsj4Kb5yHZ2UNSZPLJRmZjLpTWKjWM8zmL0yTKB/fuLqnhv2kcz
HvoleO8rGT9d4alrZLqplLAWRfaDgIdrLKE1RZLPhJCeElx3YXqTXKWkdMnW0nw4+XbhGytNG4TA
9RP9BteSlNbca4z+7FgbWUejjHBtekdlaaN7q7qex6U6GwHloUQWvYYOr0HAKicXSkToWxl1NpQD
NpLdWWgiu1IRRud1VpfH6aBU8wD4mPq8TZUxZjSPk0y1CelIWtultFNAmynada21rgu7PPY2Lyad
LEzGC1BzLYOn9uxflanrWkSFrLgerAMmcrDszFMFnuTVh5JmlXG7LStRD6OALBozH9HNhTbPJwgn
4BUhY2lHy5nNN6iRKqxDl/hLjgd4rTYapcRXRvLyrVRfpbLix0z7OnlE7Dit7NVhi/UvwIMTrjEC
DKWZb3bWjShboq3G6II8PDlOxoLDlSKRXRHoeAF9oPc2sSgdOHT8dthEveqGUHGMLmKdDwHnEN9+
Mdz3styZKPiALfsqOtXE93jJAjHMt8yFTukWCt91/GMQuQ+7IoALm3tVCVgvOuCLGFPHvz32VA3S
da58pCoVW/w0KwmRi5thRPjLOS4RfO7mLEX0CILaTK8+n2XVvvCFR/QESFfUyrX0+jSzXYK1m4n3
7iItwiDmM0ZH6x7vTY7COoccFCov0cEaRfSeew+GgXVco4NRxlseqEcoLE1yNChf2YKb0Hi7+kCV
DMt213gu+tgQh97XnfHf0DpfCKuj6ICZ94bSPnrSO24QSPAc5kDK0E0lv3MTfO+X5/BilWIMFYnL
DBooZdqVS0tASl/5EAMBZZPiBnw7L5k7sOv2/1drxYfQnaxdgvw5w+tCM3ilhqWVhUDJIAvIXrXc
A+xixf40CXI/KGYnG2/7ec1P+SayHkMYRhXy8AIXh/Ye6pOldq93KNYkDYHq24MWKaBnRyEA6frc
aAjF1U+nubPsPtnv+At91G5tVx72s+YTwwDnIKlC9ie6iFyiA6eyEz+kaswEe7YqmGsGhsaHz0A6
bGzHuuhwL++ft8Qb6ARp9eyjh4VYK6tSdBJRpHDG77a1OpVZQ3AFi9dWz7EJUxlAIKr0BvIVVzbF
jphgQLFbgrZ7gqWM/gyXP/ifxeC815AiDB+dK6gw7C1rfhAEhzHccIXI3wEc68u7TypgaV79oXJL
8cAecn8XP5OmCxbSQ8c72lWHWqEj2G2wqCZUBqoo/uWmOMBhBmqTAyOhT3EcjChirjCVheQx3GVF
5W6inxAvvTzoV6ozzSOKjvO4lbotIG11u5ee3fIE++bOxnYOtUJUOeY2SOoPUC22ftscDtJDilo1
7jop3793ODC123GVSAr1a2UyPLHZR2MNuKFDLYzLtqX9en2+lCHySql4blXPanZzNv8m+jKahthO
XxBp7CDJkpQ3DskDp8LfUCTryfUoVM9eg/7JjBNZcBg8QFAgakz2VP4x0zJxSJShnT7Mhz7Q66WV
zw5r8iTFsdteAjrLnecnUMwPmGe2pwMCYRq34usoc3O4D+GLZg6XwHLrKzBG8F/Y/u4Jd78D0Cl1
7TcghWrWNTs+v8As+ZX98YKgd2GXdIth3rAftGBqAk09vDyZJOeWGXKXHphFQG2GYStf8Fww5Cww
FYlNaaKt3aC4iOVkGPnLhAoMfteWYBbJ+kzgAHAO0zunueICMBfxaH9tLkeQ474w3jjN53Ho+OS4
S8QCOYJsj897JALi1OiysNPhGYaFb/Zx9Qk4haSqaMn2uCDeBsTF4rZ1KKdak82x/ainbnHeQtW2
DXM0fxyjnIVXOEQOHyXwZxde95SHveHPnc6SzWsFN0HG0Bdfjm5Ab4GX4GN00feBJ3JK2f7zd2fs
eKbPe1ZXve38ufL/CR3sMBJ4UzEZ0aQCzsjAgNnE0od5NxbcpYA0s0E0pg2G244CLB+uE7cxo6bD
mRKIhcWPoD8fSEaNiPA/sIZR4qUNzxObcRaKKwrFoPx3ZynisshamQP3ESo7I8qz9JBaReIFMhIo
jvJkk0DwqrSwknMb3PKri4cAsfniCHmlougIvRriDDFLF1JrxB39GwB0jUdkSDSk2FaC7Fn29gc1
ckfWk9hIMF9zNdgBYvglxZ7gvowSJhU3xcEE46rxHezzEL4Sc/y/zrTS9mwFypss6POU0g59R6x8
8B+5PEIOhMuzeDIdDmCi0Xs9A8h9N42O6y0RqIq+YgpMJpeEAABxFINGaI6I1uc/tO3UISPmixO3
23h7gqfrgniRhDqd9vdKaM2u941ccy5hAFvc+CAPu5OPO1n49SvrIZf9dIEzRGeWQfsltkbnzCt9
6pc3gtJ0AACmOjK35Zja6W4/lzTJyy/Jfkp31/F05hspsMRg7Wa9M+U7UpUZnQ1ynBmy9jq69Fp3
CFOVguA321fPCH4Ujfh8HxVGGvXdV85c+9yCjBD1m7rzzZHFBSvA3iH8cFL2Bqk+xLAY+DHud5Ef
McJxJkD7buJTEZo9bDnmQOhZDQCezlpWJ6VIyjiMQSiz/E1clX1UkJLzsZi8wV9lpAh8Jo/hyZq+
c0/BdGLzUlXjX+PSb9Vf7CoxuNfZbB2/IJyfC8KSmM//sAdRipT5QpVHNkPQJA7tMgGK+dYci+mv
h+zmdf8ZRtszq7kjPu3024OBLe5qO0RKrOm7mzLo817ks8BSv9NiDdp4CXOuLUeIj41Js87SRb78
EIB8cqR0WEGmRoz+GU+pqTHKhhlKLIhJly3346XJu1x6bI2iE6Oso1mhMeJxiGT6d72E78EY6z2V
bzldAABSwvjPCabcanzf8I7XYGVTWTRff49FsNSRPAwUChjUxYndIAOgtJ83r3Znu68BX6GecDXo
RCa1eXhyOw7adx7H9DQQ0fNDzW8Fjd3LF4hBjQ6uLve5OJCU6uivlcbPLqlIihus9MCAI5sf47yK
qncrVDHdWrisCHwVupwMrbRNc0WNVShM07dikf5bjQbK3GJ4GiEchiE61lHe0iy8abHagg16fA3X
1z3WuTAoH4hvnD2NC2UNNUHbM6/NZxOa7noJMCGBiiWzEy+JEIb0lCF1KX2uDSpNu2JP2XkDgJ1x
n2WyIdjXcQoawEE8pngoFrNusTkxVg2QMlK2Pc4dRcWLpfrK3cFhswzc+7Z0La69eyYyzjWEPhLz
uSrrlTr4Ot8htqGbXBPAec4Bm57qFnFQJFa4ihqX9j1mYg49Yow0xTqRdbBFSZ6H/hPYHXS21CwL
7+BvjYQ1paY3cZUwvJeLpVKyHiBE7K8jt9wEg1x9DqoIq+py6Rs7wEDTUOUAaXQwsKT1/WfsSdyr
lIy/KWAx2bQXC37W0NT7AmxZVLcRUM8tUp0xjEBnzKkhMhG5BZOI3COdk45GQF5D9xesMh/IFkZP
aDYO/fZoIFkTnHf0c25H5Y+us+RtmDLYYc39pYL2Zyle+2TZoNRCMos0X67qtvBECbdxZYBxEamx
42T7JZd/5ZDdnxCO3egOyPLJXL8+xu2HZqWGCzy6viCyqxvfAC4CalrZty29ALhmIgbU5I/7C0/q
8nCRDyPT4FLLR7V4zH6eIIp7ADnTKusnnULiLo8GgSMy8t6UEj93iZ1WQUlYj5Jml9lPH54ktEO4
a5X0W9gGprte375A7qDneabXqugKYW7/r8wTKZtMUJtS/bs/6RRSn/TwBIJdF5/ZxmO7FH1X/css
rQGALjF/ggVHP20Xmx/S5wSJGqGPaJG8iVZJGsvf/jAo0Ky4ZhnfwIC7MmI4hc2dqESHycBy0D/o
bJxqNZ0BQ8PcvBUY0vFIM8WxxD02aFNZXRGC60yCN1bC2XNhug0ndsIBSEvbQKDkuAaquHmZGWZG
fMjH6FEULelwpVJXGFRK6Uh+/0c8D+bmY1lKs+U3racydO1pNVPPhdbcCTq1MYPJDY60FsqGd6a8
qT4VcXtEJZT1Svr8xwF050AsE0WmDqRjgb2+aZyhOdRBBgfvHsHZjNI0b5nG7tUIejGEp+3oKrLh
FJz0tJ+jP+t71GZrMTKv/oUuzH/NQl/Xo3MWC/YOE9S3Bam5zb6FGkHD5/I/V85ba/h3FifG7zZN
/ug+VIaIZ+LEN4rluYlquqYmXuIszvsF4FxZs1RBm/lnN6bDQg9r6SZatEyZkTX6hUMGI5cnANQ0
huduFx78/8vD3PcvTREr10mzkXp377w5jxT6eVyn5Ydujty1u2hVlIcpyHBDnZqbM8BZ5bF3sufh
nKoLyloZXeup1r7n0gaGDP159oyNHFxn8mkZkmHdEXQXDej0QIqtWwarI5gmtgN0d0ERSxjGcwsE
lw4Hk92Z/t7br7SbGX/rENUq4zGFjGxTK9VAhqNi+rGSi/lWvMYBGk+ZOhg2EYdc4ljFRrmNrQiQ
ZRopT4gtzg7OdUWR6Ry9rupuSOZvM8psaeH0pTIi3yyg4Nej9sYawSP+PIzUQpdppFyj3b2a/HB0
+VstP7CH3Nv46HE6g1BWYuY1CIy5vl90A8nOf0EzMkMbaPx9Srs1XyqflwySqxTzqrGF5xaPwtN1
zqnzavu50m6Sztwdi05Pv5CGjsn/XjXB9CdYHpB7/A6P8rv1A57wu6NIm3Cyie6690VKCFEulk36
RCfWZpVFAh3wpN6uzWVK8BoyhtgEXbLzmttBMIab1dZp//vyCCEtq4sELjBNNmcLge9DwhwVqMaz
0OABlfnwBZZnbCQJrvVBh44yiPUbSVhhEuy32wMNs3d6YRdB7TvaV5LCnN+0j+js13kHnyAeqxcC
7NoTWeB5KBZ4jZbNxv09frM8nJrlPuLc5oLCZoIyUCseKI35O80bwcUKEoWw63+UHFeKe5oMnXFl
v5JSlTDi8AwWgGypjdRt25z1iqQghRfs2k9ztyW45WZKtF4AvTmIsP4Xs930nKSzCncm6q2yDqDA
wdV19EfWzRl+tNqJVC6wzI/ieQi2KtSg6zRhX/OKQLoSETFQ5EWQqolyi3LcINAUp9xw/unq2pSD
n5In0yRs9AOrfNOXwmMAMAonynnvuEB5W6kw82Pc24M3gqQYxVKqiU1KNMas4AorAuJgQFQgG2t7
VpuEA4x8iWF1RnLG2T+i1XRWmx4GmSto58tUsiM6eFawBgybs6eLrx8+E8WdXry6Tb3X5dV5iV9M
Ss6yTfqilqPkCqf/SyfOzMq7pnpsaKjl41Q6iGp447XiCGNQCxqE2PAlJ+bzuUzpTsPrST3CY+GK
iFZxBPHLoDD3R1/YSfmeRs8nwwmQCs6ZAo/oEnhVJDtUufszfRkngVT/FLovx//jgpChTlj2ZIw1
MPktOCvAAdpkQ0oISue3xLfe2kV+JD3ZSCOYu36he7M1Nk7iS94P/GsljwEXz0jyXj//Jr8KIb74
uES87gEbjuAk1Qic0mHeOpqh7w4zwQj/Nw+DtXj0deOjRT8OzJFBW1BWKVdSmAjK8KANCuRNNhg5
oS1oVSDO7GQqoGFyUpDJ1HQ3tScM8rCo01YY+2WMMY+WWHJ8cC4Mr4cawVD87qLbR1ITvHyeqAyz
O3zzOjrH+ZlG2b9KuBtWge4CsPk0Hlh7Z8Jbj6esvt66Br+z9bbvHVtz/ttHia3IIcgyWQh8xwTJ
sUekprBUNOJT4UJw8x/alVsdY13nW607vivPOCUDCP5APGDyqvzf7yJIlAfKwjrvcVfKZ1G3Nkye
jqSMMZQdvyLPzibRPOwXMkQG+Z7kbt2x/e2W6b72+75kHLsRWgmpY5WE6XjVtAJrG8QAWYefzSMn
mdcH5wzkozvoITWMscQAAHeKmuWXY3c35Y/fDA1iRXLfhaLPIqhyxmKXwSJkZJ+WNY8knPqu+7xS
SDLz40NhQP6MRtyzJZSIE1XZ33wfw7qeZ7uJ0Ixf7CdJtBHA22zByMsnRnq9LYI8QFmVMgHF0K4L
eZULaXj+qgJ+H+IFKMgjy2qGjAnUPj5lRB6soWVljz1TKKC0NjxsKJuMnKwRtsx3WvnahpcQ0oSg
Pae7t795mF4273saSa0mRSNx+k7N1QuV6dM0vvH8BU0fBr1gcx9f4Ww0pGF52E0RO4S6ZXOk+UoR
AhPunFJjiVh/+v9BPDhcvC9m7je/i2uww9H4ibEkyU3L5NDBI75ENs72ZsreBcmPDEcAw/hOyurA
mrEYSKbxXmS0j14Ycn8zT29wlcWxuwrhSzudNGDKjF5Ttiie7XRyy0krWMxFKGYbrA08UL6lYLTs
gt+k3bf+j00WY8Mbh60W+9D5JmufOGc8I/We6Ht/NpnA8nscDqcS1VMrayPXGZ0dZIuZtHPYjvrB
hQwhy4U8p0hFnOjVreq+HTu+I6YH0naWozNskhhTIrwLw31jlKXXnlXF5U5zMnbXgbICUwEbBTTG
6eR7IOKi187vKEjOt2Ub7vjoBzl3S73fThfL4pIRxabXfJK6xb/lXZPMdRjkRL+M3VaAjVxdaSz8
fKF1UCCGX8pIVnX5sVIkKtJAFVFrjI4hkI/ZDfTlCrBaZwBc1uZGQLM2uSq8PCVt40LZxO/uL79h
ynUISxb1lKeeIiT60SYTh0d7EZMbVzBLFjyj45kXsGM1ssCJ4jpEEz4T7+OFsOFe+cSIqgAAerkU
/qsS+90YEf1VfCT42ODbHPWsWu3uz1S9KqASZlVDTkl7Ux7A3fBmTyBSvThFU3AsluZMMn8KYE4A
+9mWJGTCjGLydKh6wB6apGy7JV4uOQC5CeYS3dIQgdVdJ5vyCw7sigljyVA82ZQunhbwjOGgJJ5k
9gIjkvn8KoBgLCKj1O3PE8f/E1iBTXBYbt2fnGJZHP+GeYjOFZHAXYtIP/DpBsjI68dZ6rYc0YcB
HInn78qalt9nb9O4Y+dUK+JvTFYQ5oQcBUOfD7GN2AwLZREx8eR7V2l9X2whHms1ZoYww5K7/ElI
lrHUJI2k3CpPyWibJXvskL9TJ560OTV6c6lWPNS5Xu/BLZ4uCnq+HcroJrov61IQFJ+43LbVvCup
ZjMvMG6QS1jKVL6N2klRnExDcPbRdRjLVGx4Wq4Y/Ck7dpDYS9glJmhIbTRVswvxX6ZZ1GEVZixE
Ss654NQZtLkf27aY2YFGbGJ2AGcbOR3dBdQQW1R0ve2thokH9CKFLUSF9csaCXN3q1sJh2uSCxnn
OwnHy9t1MwUgTezClNA7NXzLT/2IeoDSdNTjkJ2q36L038WX16BibaV3NMcGI6ry2e/48s6UW/uR
o1cXicPhk8nIy2hSttpb3A0PFzOvK0rDANFWhzjcbLwzH9KiQZXURIcvwhkoyTORVI+6ubZJkVMD
K4KEAAejjAUZTkAUi+V3y2GsARJlcziXEodVANf8d/HYE3VNwmUTxh+BRHp4FWaGHuM1C5OHwheZ
Kb/uVc79r8LnSz5jf8RamS2KeHc7WQAaPam2w6HDQyBjS8jxZlxTG3aPMPdf0/GjxDnwiJRNHyEG
nq028zpZ24XiNsqJ6BN0v2zsSkA7jMAPgYyIFdDCs/QO6s7Or1bzKxDvSrJ8kKcdYuF+B02MVifn
1oNsZjyVP/dAEA8IOdFb2ay89I6bn2nMmPt5LWp/7X6uAGpPnvDTsNy26DhC0O4lluVXOcsPuGW0
pp4R54PfSN+IV2Uv/Y8Nz6cpHGI8nVzT5itnyLjqwfEWr5dfoDXSvnBCi7DKl4F7XPjaW3pQCf2V
pjQwKz0vfRFfVvg3tqNvoYf2mJSOoXIDn7xMr9gkUJAHAOCcsT2ypOegfOkeGpmo6XTHt3w6ujac
ArH2SdzT6SPhQ3Lia8wtMSvb1tg2y6kr4MMpd1MeW5FyC4hG1xVN/nbEgJlOIBDq0gp/vJxtQhL5
pCftrTdLFn1UkGq8OMpOevpX5LJWqHqZ/NIqNre6D8fYLON/swKpdATXmT1+M4zYx8rtjgRfIPLl
GQMbNP5QzMG11RGo6C5MDS7JGnss7FHSTKuifkGxg39QN1gD8UVA8lfVroIeJ/g8sCuwzZUX405L
GaQuehy3MED1D9K6KN7/e8TATIvbYDhbwEmHB2yt3NUPzOUeIGlLj6wbj4CARqK2mcYgcDa6dnXi
2rXhBVIS8yvrIg2/x1wbUIdg03t4Tv/tI6PwT/NOBKk4m5BLKzOe4Im7jYIv55rwY52YMDPBENox
MKAEqwXlGnIn5U8MN1rDyYJmIQLg6NkR6BMvRj3M1N7z3tqNiRrhohj0NEUjZ1jp5DvlvSWgsV4k
AJnhaotOZr3TvzeDyuXtTBdDqfpFeFYEtUiavkuiKzIlXuSI3XQMzbBTvcpLu1Wgj1q5qxIuNiEk
GKh9blHdZ3zk3DzAwT93rrrzmZU/1YFg2/BoPL8FMsm6hUvFPZmUqSR7E3H0jTemrRTcsEHd+QS8
oaFfpQ4kS5Hwkbt+SUi59Mank6fHXC5iVSVEdmT67zki2ck8Y/4MSUN3EKHUJ68XRfAxwAivQLBK
6H+pnQuiic8TupV/JsuLnipydH/zJMaZQGtSJZFNa6JJlkn/V3neJOc/v9yHr9PIqp8vbo7hLGb5
DCpNpMkv7XQ0hjbSvgHAwhtPrlsJkJ9LLTdRrDFe+tV5cUVp5hGNoj/F3GkoAkxB5x2PtfvoVy0t
VYMLTsQO3yB76wg82IBKWCAM4LujFrvyHRKgoeD/HAnxbO2/W/204KeyDd/n+5IPCKqs2+gTglLh
82IAChkX4JSWsTise4CxEu3NVDbZfXR0wcGsSEtD2atPUxDKNXYHITE4iFJ1ssXJWKkysmQ/lzsX
OogiIkACn9z8egHLUyDlnQVYo6xYjpGBNUZwyRhER1sKS7kbzC4MrEuaqIbFfcyfTgkBehule/tA
dUp+p/CmWrHqUTrxL4/DAv93FIl19+m2A/xwJP83t9U45/z6a4XxZenVK4j+q9/hN9mlP4KUXL76
yzMoXRo0Vjh40mj8RUtfBoMcKKnKbWIAiyU++uZedfkQnpwkJfB5JYVpM+ICFsnlpfmtOrLZcyWJ
SKlzY/DPVa9neO7EbZBcKQc/MHAmgmbQfa88fCUgnvcumUssoottU0sMdBgM0tCxqsF5Wt+aulVL
A3WKKN9x0BJpvXQhtOVpCK1f9BefzSWDiRiUAh1mlXNz7vHT24nnt/ScKfAzvPQVVUZhLNnCZwpq
qakjLptALMzToqE2oqErcvIokeITNNcXOUr7QVUHaEEfBkOhqoMVoMaToUUPelNmv1k0WndSCDa6
eVRTS33K993XiJBVDOlAhw/ruDGy+5E5yMGimzRcbaStOSnqQKFFFSSp1fRz/qNSQTioxK7DrTJq
gZp5oTgtg/TbmLSDwjn4Wm+DZss38vFSlLWgPt4Ory6qc6uM3IrzKfY8QlFtW1mZ95we9Sst0dE5
9Lp96ijQRwAHRo41IMDBRRVM1Nn9kpVJ2u7qtde+Ehv9zfF3HlgStGkgwhlmdQ8cT8X68nAkDuoX
Sm6vC02pUzgkTFJxKBcWPTodYnGaLpLkIjpHYH1rFHNqYV3MmGSa1QvhVP8+H/aFnxp7Eqe+/SiQ
Qno9LFEg61TZvh0QbXFJls89rWq0gY+mcQkfNjh0c2TD6crHE/b9rsLrH920UZ3ZH9bSxcejnGV/
br8e4Wa6SfYQ25J+Vcyc3ukIxWhF8UpcbddKVPDWpHAy4dVDnW5NPP+xMnfaffrqBKrqjdI1pr90
plWLXHgJqgxcr/iWV172Te/f7olQNLBvpXFxBiVNGLTK82c0oJ4p/FrhCJ5lTGbl7L09jg6Q8QVg
SDe7ly/Dg6Ld03xWh/c3wqFFr1YaVL2KSpWgIearGJL1RK3vUG/Jt7AfxNAaSHT2IEgx92gCmGHD
PMgWBR0FJWQaOCEiM814WEnvy2XSVrmihMqCBcgvUS5GM5oWNtXhUMAuZjsXtpMmReGG+SFP3EGt
dJxbRLSKTn6h/mKr816LBupcBoxD7DHBhUuZmPY9JG/4QjXtgd5WR/53+TY6VFTHdq95wi1U6bs/
oypHpKcjD+YU1aJJ78+3mSrSxdJfvn6jHltZUd7GEg/IDg0rei8mh9JkKRvzgEMqMqkceBfQHrZR
jbf8zI1wQmApt3FMysuaR77d7NHp89rWzMKePZ28NQa8DTWLbr+OjtfVCwGFR3gfE2mKYwxpOvka
giEClp9mtYAjk+ebXD26nY0rYxnrYwt72EAvyw5HYziDoQURi2X+CqTrwFTSQpqpsvu5UBM9+O5R
13KZEUtohYDD5jujd8yn2T/yKlXaqL7HX0U5ncmaQDGzoiPjMmQam/EZIGtUpzsAOBQyYSPritHV
4qBA+U5a/zZNjnMtznygfn+8CApU1f2Eeg2+iEu6Pb32uBjLjP/0cefKz/slSQ+AJ5CMFC2Qnhsq
ZaNhcwU4y4IBll7EzaXo2CoSrYEESZph4hoq7Cgi9jwyoTBq1qkwfRcHBJlCJEwYSQX5FuWZ/XUl
pMiHQeMpz60n25y+Qfe9qI8NufVHzWJDp5ANUE3CuoOUZrI+khWW/vZ4IjKUPS7nbZ6FXa+4hAY3
Z/5dDSzEcO34G4+30VXf7tUaTglM2rDFCGIDsxQfYVuWejwuNES65puHNGLv/KkEY9Rgg9THufu7
Cm6uo9EqUTYpYpL88iwygfWYd6ZCickONPBEuE4iw/rIPdiVKgs09BNDIMpPVc4+mF0eeSlwX9+C
hRHkCi0QnYH8Gj3PuwMkEg4DHy3MZ0zwmqakxEs1vvSuVXbZhFhhBKGQFNIyyFT4zG8PSTYUA9iH
d5ztVqqR8Pu5WXJjr0SoC/yh+qIb9uQ2TVW6/8glnkCup5ePCGL5KAziGmKWN/7lcFUuRjuIDUjl
H/lgv3dzBfDmu3k7nx6wAwN7Qv+xP37wx17XOYCyEJhDwzDGv6gY5Q0cMj2vbg/VAP3j8JBFgJPD
BThcmo9Z8luZ/qfHNY5nrINbENrwO7gMiKky4Fe6dVBOjP+pVaq9Y7dsQo9OTzevHYbhlkO/LXhc
KjygeMVjmwIxeZV/I+9a9VJoWRbDqvPwnma4hDHwJeUN4j/Snf+cIbRQp6aE9XYIju91jMPMnUwh
iXvXHcZKkgbYMFNS8GaZMfJ8NSPnNFbZ0K7gYAS32H8j3jVaBwC6IVGtr06pe34MmCV8YpyeOb2+
UIvLqz+lo8eyHdRQP4piq20R/Xku223Z7mkr/LIEoufcThjYjW0OnEBaz7ShGyfrkYnebq5wrUcZ
qplDum9p4wRscuYidnrA10FUkGaAoW6l31CelPPQAsyuc3M3T1Ui29cIexeDCXSyw+l9GcgPC7nL
NR49tBjTFwgbeRItH+7cn384SqJ1QC/6oMdvV3E9X7k+WNRyBoHVbpO4smhVazyoa4bz2Y6REXcR
WtNORqYb+FonleDsA9Lq3Fl7RyBadt2epmej0Ml8//k4FXrmiP14zg8R8S3Fie7RUiMcatIgJx/u
nS85NALlPBFu9oqnPI/rbOiAj3OEsQurWjPrp9EP/vBZMmQrsHhXuICDAabwu3h+OU/DfMUYLzUl
d+PXnN9aQzoVEzhmuQ/t7ijtD6UHg7Mo2UAsuZxInnlFP0LIBP3160G/OaYt0yg3ghvErV587W+U
uMLXcyZRd7xyyfgDgqJHDRUX0DdYytzbSn/vGzZTAWjNGWv+S1aXmYrczo9vSmJE5DZY8O5culaQ
At4V3MIY55k7FgsOLCgl2ZTDm7Vg08aMmGVKbt0ZDRcxCOSauXgVlJlcvagupl0HOVycxh5km0+h
6xODuDjTYd4axquOQCzDpEADFtFD3tsdnvWdNXzG6BVMJX5vYf/eLW8bI8FLgjO8ahvxq/usCUky
LGTWKaKBuuJDn7yIxApw2M2NEoexWdM1aL0+H2TYEhlAFzpm7RG5/HHnwDzCjCFAUC247wFrF7Hw
hYAVXUuWOG98YT6/3IjD6zNIP0ik5Dyq3ZLouZ6UDy38EeZDwTDdA8KFDEAvQnCN9IaPatogcaHF
6UJLA5ejaKP+NbuulAuWyyj24h4Vtxf0XzD6kCwzu0hXNqMc9rbL8uD9VWr96jv6zFtJdi6Wvu0h
RALrMZwEK8J6q0qVerUYY/ztQcDQ6YApzhdHt63hSQT/K8JBPTrkdTJNThDHUby/1XV3SrPbtPuS
3V0MDBjksCPsjzFl7qVcZbazBJrfa+m0MFt/LLdKSH1+yqXCs8j4YMyAh5qxODznvY0zbhvvmTfv
ypatBx35KcmwEprDIU+Da7Os9mBO0OzC4861wBIMbf496sgTS3+/0gKpsci/4nGJpv1467y37PmM
zcKI1njf6W/wmwMmU7rPJ1dWZpyxTg90wi7OJ3QJtMJFxjDTeIfhpTun3GSOIQhlnFByRdPikvkm
0QuEPqK8x+oQIKyouqn6C3oHWqr0TuWHUxGeuz3hxZRX6qHE7/pb4oLrBTKROQjGONkqhIsNf/w2
JLZAOfHOpjAAA2hWXfq5lYO4mUC3ZVsukHxnCS+V3LCbIMxxkcvcdEyny64JtDlGOXeN0G5Zxnet
Twtw5hZrITZ/wVmhh2/2x47gmk0QthfvH9gQVqeDJSYaIbfnQ+7q/XpB13zWrirhpEWu07pM8T+M
yDH/Dgr65qnRoYuRjoG88wss2Xkr4lHOO7OI08PQgbr4CZSuS7l70g/9vh85k+1aXOojw6E/ogob
5cygDbXhcDz2VEfvx0Due9eskQtT0rCd1q3Vcrk6AHWj3H+Cq03NJWSdDW/yzXiG8yqghSNUn+pm
9X+BSQFarm0zoMY8whuVIJluotOQK/VEEySoHPwyhRBCY6PdIQoZ4ZoYhNAbB6ER9B78CUxfVDwM
qL6DY+7ntpkE2PD+4pPs79nCfrw47HxDFloQ4EidmCokaGL9CR0ZSSjwLvoBvU+tlEs+g8xgfk5G
UKlHy9X2Xy7IKSD8z+YCHoIgxVZOHoklEE8WG0PBg6IXpaBs4Sky1H5jYbQ53BXVWVjcFTfcbB98
90Le4p5lhGv14k5NxwjLl1HRQc0Rmvq0NJfFI3o8/RdiskEiZiiQfUqxjiGSvffZQ/1SlyJKsUO9
mYPJGQYuObWpy6D/ncDNI8s3stbHruQmK7RYxZ42SQvUhPUkGkG+LuYXBK8+erhzMFLf2YDY0zAa
nDE25qPWV54GyOWzpMvurMo0tLvXoZWS4ciaz+48tRBSElXYlgwv0tXx6emS+gPfyelkY3ibVima
YS1/AuLsiAlVoRCQkKZNUX64lhz9WkGX6WlyJXiiNYFEkMAYzI7yoXITNGJem3FkZuqiVm5U1vwm
XDJL1qdFhfYqiQ3Y1/2UjbQ6ncIoVIK9SI40nJFQsfA5umPtMTHsUuX0/N7NXZx38+0G29wnMg4O
2fZPc8B9JMKQXH2fq7NoMnSgzCK3ug25lhLifarSDpvZiaWub+J5ja2NMFdLAf4+L6L5KGmBPAby
EmGNrs0yRLwhFk5kAbFhmHtTM9xqca1fqaTvwiDXPBK3mjX6Bmdzc+5Hxwnf3r/G7XneOSqBVElS
Jv3NnFadH+yup0rOZFTdQeJzRlMc19XGdvYF+CYh0T//0XvGeF4lSJko/bCffqrRYKtoE4TBk/pz
X8V/acyZfa+vt/YHsLmxvPQ+WydshL7aLVP8HJixOOTczUxYBx9LawtzouEY7X+X/xzRGJJI44pS
Lgz0zewBisRBhy8HcytPYuWxsLVOHJ5zZ4ki/Q6kVN0yWAv+smc2hQ+/dGGyxDa++rdtj5WYXEg7
KJICr1fcVzUXO1BAFAl0k6GWCbyPfRpq966UFsfom5mOJozUoDv//LO3r3QxvsE5X4dfaLecE0Iu
t3UNx0bJilYS4XVyS0rjwlX7/cscjLQQ+YB7pMbgiQ0HzwDlCiAtte4VwoC0kmNBILH+gumLmGzk
BWlU3x/V9tGHMZI3UD9IqseEkvJ4H45drbZuDzzhteBf5wcJFC/sY2X0FafpHfX/FcZvGwAdEocz
dK9Fv03WSDb5dX9zLsATWY/3LvsXYjzjdbH9PQA6H5nOCnfwufq0ZLzCKuXRicr08qQC4LCsVYHs
4JFJrxZVO9GS49amuDcaVieR+14lQwmxDxowCVD/GTwe1YuAE9/1pBz3Nqk37dbOFtvws4q8vQGC
D4qodJipssIg5qzRnSu7ElHRcWnob0L5vMfFHRq63zjjZgkmhDN+bX1GSMlYNzaJ///bcj7D+t1J
KCji4Z8z1uoa4sFgETCj3hYxi7GBKdWsmAg53AILWRoA7GQ/00Y0zIfozstww2J/2/PTlDMTcU3j
Naf/nQWgW40aQpO3osJWrfAbq6HGftFUIHI4rrJABQeK7qEvUThJbF7Nb1FGelZsjptOi0CnxvbC
fG7K/EqN5MtJVPtd0rEvKacZS5KlFO05pfOxcQuQypT2VHo87ecNNb4lWZhffDoY9M97J6UIuDVt
LVOKfzZ/X6K1yjzmRqi/iKt7viN04O7PvguLNt+BczLNyhLQrFsfNYbdc2eQM78RfleJzRthdHdy
aP0AZP9WUaONmpXNMSpk7gzm/Thz2TI8u8VaUAR8h5hxY5BbNHIjgRsvw4/h+3q64vsBXrhA6dEX
6HABDFPN4YCVb9EwPYghvLEE9Jx4y3fVltbs4rWMNCBFsq3obQUCTMUfbbKhJtZtNUBgfTj1qKI9
pdohDh4CjXNB27Urdc9QA9XGC5V1RITQlfpryeAigNOYHL3Ll0h717mvYQMPmdJG2h4bKbEdXGbS
UQUZqZ5TXtpvWyQ4sZhPfkhezfP7r6xfJqrrLSUTtMfY/pPLf9IEqdrEccJmOSBFuWKckilLI5vH
NUely6amsoSObk65R3G3XIlDk92tWuDByMg8EAbFeiTcOa8IOXBQLq3tWhVvt22J2POXscLx4bkB
Jli6b6lAlw3/yKwXaWrgRD4zN2xGvGVR4QdjQa0PXthjUzFEN+2pocZkS+bT/ScJ2NWWC5yGyeHM
qsf8vCsHkQIPXY9w7r0g4JQy4Nb0gGU28C5Rv2wGOcjM6cm1pGXUMyfiB8l4IuaINlstJdDZbt0q
CkYvNrqFgJ0ch8bUQhnD/DM5rhc5E6yqfRCso2AlwrVDptUHbXzqG4oUi1GPzr5G60kCbN6bshzq
LBvdl0IrHvu9xLhPI85lUHeBpKtsn7VHJfxfT4dIXvCUre15wJjG4lud/bhFujbZIdAQVwihBQlm
/yeZ1vTzeEEKE3G9GBYXPsDCiobgCuQwD/mNyFQWIjuxqjwi6uQYd+8NMRz5SVgoAcYpQBQwlGWT
wv/7xsp7YIcuAtOYnLVO/FBhpbo4sNv3wCiP5KRa77v+KSZrsQU22yGm5dcVLvR+X/5B5XR7rAbz
hc6U2coS8g+1aJXoKUdKOKYSXamw1WtYsxPVm2LX3P2Oq37EfEVFFrJG4MiIZjczQGUeYQqbn2g7
XqUafp0YprvZvxDfnMZk/ZfvYjCdJoJj9v/VZAGSYpRsSuKCG+H+kiQw+ECwW94nzccC3T6QbNt9
qQGx9PQUOpTTvvptoJxlhUY8XnPbmOgqyblQ9DcUI3sQBr2uuz8Rnz6ovJltZgIqfTvqCxnH8Bv+
7Qf5iVfJelUapOhXCwXolAqkiab7utlyC4VXeSKDBBcOiSuu5YapSCj5yxGdpF7+2SnfSwqA4fmn
/gEwbvuVKBAkklkNhCNIF9Wx5YRd5jQoE9Mye4y1Y05Pi/BH92Xi9UVALqHTgtnme/awRdzI/v7L
i2p+sxC/gbQ719z+yUAa4DvKKjaKjIOK5XZZIcii6dLcHJRqktT62xZaUs8NZW4ssX+d56vkCLoA
U7F1EYcwjdVhLCerDpCUwodnYTorAplHHaYRrYPdVe2d+Vrhy8dLHXz2EQzhE+0hvkACm0AiC9yD
HOgqmqiflAUsts6WDMUq/odm3b1w57bJn9o1L9+VbRvNw75rWd5U5UkjBRrmHhQ4J+2Xo9lSdzsX
+v5pf6CfH+CvQQFUkhQKj47wQTuQh3BuAWSFzQ41pGcjgJg93pBay3bkmIMfQZmPuqkpjallYlhX
eGCTKFvOcZd9ppCea2TJ0sVo11G9f5kqiurJOSWSvOD7U4SCd4xQiPH1j34/57+WlwpE16+pFkfE
z/Lj6qA4gkUVdpZUgD8vTqiU3JUpUWb/91c+mcjw8mZPkWGuVrGPSBX2P6E+2ME3jVfi5xajH6aH
/Dwy1+qV4LVW58R9Gz26npNM+phmTLtBsLcfuA0q7asrRU9nix82gUv7w40uT4/sAhPe4NmTYkaq
bFfvb8HxiOztryFW+uSDkBoEOq212r4jqQsFrT0Ugn1pXeRb95GdKtGzSGph10tstuJyvH48W79m
Tu6Ou8K6f0Ebee5hsv3hQZwPKtY/z9IN3d7VEUi24c8XEbYd9Vsz4+l1QrFIIAQucmK5arqB4mJe
6qp1eVFDiBb0S3WBTZFuHyJwBRXE1TCln8c9ICaaA/lyeaJFrtWW+KfRt9hMCfkt4fXuIzqk++Wd
B2KvaQxndV7jCLpCeagduNuzjzzIWUqL8sNnLv3+8KJyP8O5kqdpvllqCAsqrQcgW4JlPkS0pDAm
oqcDdZm2FelEfb+SJydX1R0xwivQGW5bSHAxB27wKCAK7CtltcblCojCG2/CxjiFw4YW+16fYL6A
4m0GY73bbipNIq3ty2GG+gEpcJAbA42g2X9IsWXosb9RT9wqtR6Mdj4JWYBZO6+5mxiShYpCm9DJ
WlrfG3Jz/e4kervMSubLIEFebUFxp8vGkCBkoKqNfHhjaRe3/g0VNnvx82ZXFetgvSyyVVnfBKL0
CCIFxrU/7siusbreK9+DZGNCvXSRrteAXiog1Y39Pjr8VwmwCbcEZBWkB/+RUqOWh6bvkIMPyDFk
NgXlR6P4cEtEk16AwllF/iXo/ScZVYsggUh64gX/W/jLkb6SD3N6zzbqbvcsW/Jxs0+eykMqmgwm
5Udk/ev1TsPw+Uj38Zoph/NIu77c2vfait2H5ne3jPXXBGdPoKvEmxIFFa6myYM3tGpWoTnC0ZR7
qYU2vNVOf0/rEjnc/cIoJjvQnZOTfUrPysISet+AOVJtJLLVf913yWAgB2hjRC6Im52P2U/h0+pb
TmqSzTrLctK1rpRnYgDot+7HCZzx63b6zAcnBsLXZRmxsqGhQm9v3wWBvh9Roo4OSjSjnhS0IZC4
u2D471ZXuq1sz9+z97XlAqb2EmdJFhZ1X9fbjo4+lXm8S20UtT0iYFXjlvcLnOfB0RiM95EFZLVw
1YAEVAlrF0Ufd2NweWRb6O6Xquhf+EM2RT9BJNREM6/kE1S3yXiI5JhsgToDRVCGZnZwBJd0Mz92
MVIzZfty8EXLsk3HIdatBsB9OFKk6NhzX6pTrTs6XJA8MtxPlc92vCDm6WDzPIxtt8NzCuIGm8EN
DWmf+VsqSPTWrgXoH09XL2j5FTunqxP9WaIB3wQzUIhB/AN+zi1t1r+wEhCcezcHY5dd8E5AmMD8
2Cvdc7LNNY+CdjR8NNX4+7jW8/vQa92VtxI13Q4tayegdaX9x74+Q0oByXvrD3TiyZkmlaV/mnvX
15iARzywZq87ZnAuCjxxBZpgkjuxhbT45aixrWDvNRswzq+btyR7VfVnkIqPKYLUEZo9UeKJxidr
V7ddFL84TArBDHVs7Dqs6ryMwVPQbP5p2lqcjr1rf15IikVEmkstO4Nb9uYTiMXFvmiJR29Ope4a
hoEu0wr858lFSPigQeNNHxBOoBFSvKEP8OsbUel74IOFjmoawzMqPonC1WKo/xR2rdwwln3HV5/X
FN9TQbgFORlHb36tkDxKvsX7xEFFHJBVCb+KzA9hOyiibsSTsu758EARC7CacwdkfZXGY3j+vYtt
hSD+belKJP52v6CnUUWXKR3DFzE28ebpxGGClhUnB+bBBuKk/v+G+8p8CPU+G/TJ1w27bZ/CphWu
3UBTu2RCU1TsYLRwsDsqNYzT6aoJ9zGfmvTp4Ss2bNUCYNPaXOTSqLEL3rT2z7Ajo2U7hkmVsLLq
Xz8nbwKV+dfXwQtPNJ6tdvqEoTUz1CveNfLHcWSaWkZJ6xDcdSJkbQo8rCDeIx3SKf1fomCOQCmH
Srpn0SCz9HJXO4HqZ/uAuIod0cLj9UVGFGv2mk1Q0w/n6rACK+MllMVYkrcQAE0QPBHjkWZ06lHG
yeVhohclhDel6FmQs2pqHShB0AKFfC3gm4M0jgM5FVx0lNRbouei0oANsciXfuGE7Ys95uuD4EPh
RzWaT2rd19jFlLtJs55X9N68Xt5kSwu/ZkRo1/ncqht+ZIaGLGxJhYsv/x4kmOP1t+bBzMRaR0l1
PTKCTdtWymXYsZYKBlajh068bPWyYbCKysHTRk/G53R0HKc2raiDNkKtaPfjmp7KJSxZdRaCQrAQ
5OmyXF1Op+zyWlfeQ+Vw5p4d9sq40JZZr4iifdw238Wt+S72ONhyTYjkIzJJaVWUq/ejd7fRw4VE
JUfrpzcQL98NoUlbzqN7k/Ml+oAfk6En07sKQzQYYbqgYMbmFkL24bodAiMT5kGfw0flQ5iq+Gbv
eEeEWsAB0arDuhiOS/fwQPp+IoOLI7HmYKVI4zkOhJo5jxQtRsNWgcqUJcY1v1qPY8yY0pSV9Ch4
uvLalePnFJZ22eKRwDXvd6e9xupe/CJe/RYxq/ea0b9In/+JQiLnaZj66wZbeKNsMOjXVD22XPi9
1vgrgAu9munsoY+Gvbezxm3YQqawvp35Pf/eUDxquUeHby4M2sZNHnTJcsWrDOIIElRKyjwaDAaf
QfNH+WEgfV+RB1WcR76SI89FnV0lRLtp4lvxaAbDYQpqVG1/W6NOaYvqEBCF500L2+T5v2KZ/FcH
EiQ1etReqD800tIchzIpNjkHWzElcHock1zQxYiShQdkrWYREHkS8ITpZAcF7WIEekIuTIcu++rb
Gf4NXLs4Ube89dpYYLogN4hKGLRQuuht/nCjChuTDwIrX1VgTfm1McYTdnOda+hHiqfyGvTeywOL
3oc20/6eoiBXiYOnXPMjW/xOC1Lq5bZlcmuzmyKovR4UdTEG4CT4fxaINsWE9ac2L8JQX6gF9XK7
LBfXRYDF6OyjxiM2YD6MnvQ1uUT6nHSwsmCDVaB6D/SuXO9vaY2wKfur9SrXDOolTVJC3X0F505W
2XKhHlaGNfvj8XL7SBF/bvV7ler+2jWm8PynmoboIjj9Wxo1vYJW2Am+fgny2k7j4hZr0SrAMu6G
OKy60Iz+S6916d5NfzvNZpkXretje8q9WCmqPBIJ0IxiSviNmjklnDSHA5FBHHndh3AwbdZY2Da2
78ioFX4HTeG0JnXAykJwiK0IbnDfF+eCPWkMguNWv9b7pRKGvUynkh/YuQUvUqQuurYWelAzZRgi
CXGrUFbvBxC9AvTKRj7vSS+36kMFvkbTfWf9r3UyuJLElmWrDGqb5tZn0Rm9bK1PKcyz4RwVNZQt
NaJ3b+yBTLBUoviR7KGdPpojDYzuzqwBcUfTmGZH+r7oCXX0tuu/LHRKWg20xRVjRuL/qwao8uvf
Stxd6iY1lTI8ElqIxUrf+1ZZPgbdSab+SjKYvHjHMP296CVD1havZ+syE8lRirJDZWXnyxNztbsl
7UVp5WkVUq3SQP81TqFl63bI34cntgqDBYTWmG3ks1pclkBM4hrIcrfdLQuBfYQZCsXw+GDH1Sq4
MQGZXkaSXmRVYGY77m+57YBcUSMqGD1SDtq+k5JxXXwttFAvGlYcOmF7w6bJJ73RrXNWVovC63uf
tpSI69XcolN8s5QjUhN2sFK4LK4G5jk44gbONfOGtxKQd+AFtuYLPABDYsedtDDVMK8kQ0HzrmTp
ImQ+oqkF7zGRypYvJf0QseVptqc02TW5WMJCVuY/18smavTJwfGUCORyZkiglG8PruauE0R2iCeh
D99wIP0fQ26S0JFohWgHfNDAfPIljFsDFA7KC0QGGsPWFsW4vs2dG2YllbnwXLeq75V12wOcQKJ5
EeOro5Iyd/TPCUz4EKfd2qzoaXABJFqRFOFnfXRJptp4omlQ5oNJEJiDRvYLhUp99uH9MK10ra6/
6KNYrHu+9BTJfXI0a+mt+kjjyyzVU5J8cRslQb/HBc+UWX03cB43IO5lNMP3l1tKKWC/XsmgZ2ob
68pWDaInhOy2cO9UNvoiwk47LRSK5snwMcAsDN/JCcoXc06TWVHXLDTRQTWZVwiAewb5mXzWUIc0
Qs+TrLPfz8/30tnbCMeF6aHe+yMhxlFu1pQ7pVS3KJHGShWSq28BjJK1lxtNHu5kREQYJKTbLpZT
yh8VMrXgzvJ2GXwxLaH20LLNWJnGEEHyKLSYqq1CaRMyQ/v1DA3l3u5NxepEOKmRswRrjJF6KTkC
NlZHpU2pQhY0O/2AeHNMm2uJ3EsIfvG1Ec4qqx5qVdN/G8b+/THtM6BC7lEpgsm4tlIgXihP8anP
YFbbAoo4O1ATl7MY21HBjkLmkw63wP54/zPVERDK2WhLE8kDr5SQHLchm+aVVS9rZV2dDJA4L2kT
9c+rskxf/D2RGslXJXXp+GS6hgAPr292vTwECuv4hdrj6NcGL52PDf0RM81s0UzAlhfYifls0+S0
NuloU0hrEwLV4n7kwIP/JLbp6J3epmuR0iXWHW2KdaAVDD8CHpmfdYmLpshfoE7pfQjbZXcmi9sX
BnJvueai6eTP5ZXnfN3nPhruRmRViHuOmWRFSzLS5GqdJ7IOBERbm5LURJNwolhhR4rcLbekKpzh
/jE3MBaihbCTQ3BSKpU3KjrCHgtbNOiZ4QuGpboGb/Eq252Se3mLSJuIbUe2qSTI/gfm5FFTrTq8
i9gz0cgbDvGG6rdblF1vP+lYxB+XI5pz2QUrm3/Gf3Tt8EFMikTFwbgAcYitBsQ23KH5qZp1KwUJ
nzOt60rO+N8FA6wpwflfiDmkfSNB+hGdLfQzaDOYdr2Ocpiz8hO51LcwPz2S8rrg+ATASbkj/z1O
WPuSLDbRH0y6OwEKWY50e/b7zFW0DcU3N67dQyqiJ58jQ/5DKburapDpABjVCnk94fRYkDMMoLLT
ef4plxn5WBJFIuAlFDIjWMW+7xVudCxO5rAHFZVtOfRRMJhy1fco9ZBV6iQbUDEU6vgx8f5qQWyp
E8PrucS4zGMl9wN1oMlZy2OFlJzyD6psNuDVDU/Vk1uJTnfUFoDMk4nyDtevNTFsLYXG9foLwvu4
JhcCrCbY9UqROxbG0KYKuqn0TxveU3oTXUYpTvwfRN8mJZgjL6ste4qRmZjMVDerEgID2klq94WP
cIBXAO3+415X/OTgaUEzgylb5Yj4DCsHWXkx+vUtYh8vy7R5/i9ao7d/jc5WQGn5Gr3ZHt61JXwb
cZ6rpfT7cnOygaRH0zzFl2AZHgaiyfvwEikOia+/IGFV+X4cC3tnez//AUyqoa1dzFE8l8zv3dJr
Mw67uVTTcbLkWIN2uZFGl5W+fwc4uMhIhLLJI5gzCc0WwODcfYuGhAzKjXNpIsKks1EY5SIwELQk
I8Aq2VyrtlVptZ/65aZV1HOw9Y2NwFzcGYVTaeqO5no2z4V2kI0xq8pT5vDXZ2XhN5q1E86F6xRj
3I/O/AXEJSJfKU+4byNVASZ66nreh4OTWp3WGEsqeW45U+k0636BRH3jt2hty/EJvI8TXaJ9gAuH
JikNf2OlaSL2gL2woxeMZI1JI1Tw/muaE+HmX+uZnQfMGsa9hYT//f/cCK0NTUbQiDee3HruucUR
tmeV5gsGvhtEOijrANpRtUVUcfYF0IlfxMdj7XgxRQZ+NgkzxwuHGJOs1krUzCrx3Xibo+JW91B2
h1JPK8yLxYeeI/uCK4qfZ0Ee7vmNcoybv8ZuAA/yhanMtBqESfXRqUSRsfGXsLPskX7NkEkG/FuH
A5lrAfboFeOOTnfMioSgtbQR33OOSBsnTqbUQWtsay0Q2HM+Pge/tXe6Xa1YFbqcUp9V7yWxR2GR
97NqtcSoJs0oAXRh1+MDOgTG9kneH+/cpUBbU3Bi6pDiYRUWgtBiMCw2MTxcBfYo2VD/v+bqhXGE
bRq42uV/OYtlkV8RajN5heN6qA/KFSWpsuYMcT3cMncwMsRD4FWymm1t3ePudgjhsl/jwxcCOkin
xMceQE2xdT048hPdzoHPHj/6hrEHqYhWd7KbWzyAbbAKwy1NSpOHoTrFreZa5EAPpUAtMthNHbdo
lr89/2hnUwUrEoqh+DK9VJr5/dUBW1meL3x+qx0F9ovwgkUBBVRapcZ8uWLsoDHcgGpv25GPd7VJ
46MRw2BTux/ZIrcdebWx1wiycSm13DsPK+gWxErq99OtxDUniYGDd0fgU2QjzUUBFXXqbQF/knx1
ii+jC3vwXPFb+mI1wmuiYt6ZvhDHu+j96T9IYqFeYJAHFY7+eexJokIzXt/B95yZbI3jlN9ZRydb
UN9hZ8CT597bUZgOfl7J0UtKLjBs0EKkRdgnz71Ulec+fW2xy0e8852frICcMul4QyUiOdG1sQp6
722b33P8ykbTmV66vTgZCONvecjltGaIYH/QvbV+lhfsyVLH4Bvd26D83p0oxmrMe3lvywGvykQY
5Ddko06bHyvqfDS9rZHYROhEJ6A0cXhHV8kyfmjndZYQDMtoPrfLtqP/619d1aZC6dIQIqYcNyB5
sAgsGCHnpOYIMcUb3/HE6gsBv6VqbRWrIRo3dyEh5rgeS/eRPlgqkEms39dW49Ai+APM4+aXSe09
4yTU71gpWwNsz2ktwJFb+2t9O8NV874D9aqWS3O7BpSvDjv6TfzUb9catwMQ+Qn593YMeyAR6ZaQ
Ut6rEmNoBxGFrmV2cwo08e3NZZ9pNIOer0s7nougd2a+/EfisOJWX0rn7bgs3tu2BLNYIfwKbYan
Ng9VG3h4Kw/4ZYVfFYXZCnlnwXm451CfKFr3TYILrGy2mf+jJRKcrh59DfQitr0qZVdq3czbzK5f
H6dCtN2TTMh+xctqvsw/xRnKKYBR3naQVLy9oFKICeZqyA+o2BjgHdswFru/vCPUOpcYxbvxI11D
phOpSHd0aeoZf99HhSCxTmfCYFYrjWHlV/1QyMl2kbUzVBfmT/r6ZFlWCJMMxo/65bt0HxgpGoNl
8hoxkHZraiQx7j3efl5rZn16KTpM2+9nzh23P1Ws4qn/Hu53yc8YU0Vn8fph1Y7+MeyT+rs7pfxY
vh3G4x8pKG22GWrKtHpmAjnc0uRDdvthVwI/+3bytx1s8aAeflowDwS8RU3C4QBNGNXvny5kwbQs
gJQSj7gDe7NHhituOgOFcJGlAxXvUv/xAON+Q4Fr9cw5C3tPXdk0QoCEF2zxB2uwJ9ttMRL4QsS/
SD5tjfnX53KBQuJLiLjoBmXK+pRxkCVnKbw/O6uFbcH6/gLIw+PNVkj4v1EWvDvQBE9bH7K1AzU5
NOnA5n7faokYpwqqpC4uQ5tTy31ib5z8JjdLq0kQ6CcGZW7bjtMjrrZcscVRUoCEz0H7vPY/mrbG
czAT+nCub5NSdya7jzeuRrC0dwVlnqTEWpHbBYBIHY4MGzW4iJnrUug6gb+PaGzcVci3nGiiFLzt
sNi/cW5/KdYRRGf28K9ubvm+OtjkZLOZSXBLUqFKU5gbsAg2eEuM7HAjur78CXhkYr9hGPszSSlG
z09Et14gaIFUxC6PhztKKyEcy2o43woxnc3jFymoU2d7ygmwzK4mLo+cwFFucLNMQrwj7DBfTsvj
jayy6bfSo1NS7TzuEJuPBM4YTHYEUxiowHWHqiqTVQEaFd1XIVnQ/PruyvxDRcuq4AqnaIkSZ/oB
oAIXQ3FjVNjd+lk9hLwZFGYMeltGbcafQ2oYgBQ8slhLkgMmHZXxLYf/crOwjZrhyEjyY+5BTRH0
EThqjyEcSfTU7+NLi5ZBZQb2Wwy5V1RvVNo+QzdO72VYPY4LodMoWDXHjG6AqR19YDPSS2Y5kNYJ
nyFcfjfP1iEnOUlKHaMRpXT39fxmrw0LbMSgEqPRVG5msEnZ0m4gf+NneQbyh4n2gqaJEtMpDb00
d1s4SoYh2rRx3kSYDeLLO41U5eqng9ZHpWkpinnnjklHpDf9tmkdKnOkU+Rji4oyzLYGmgNj3yHq
5DM4lVE+09NFT3rClbPrylAPjvDdDNeMxx/ZKUPs7eKkFqpeKRchlyjOJNMrAB3m5oIk8k52B+Yg
TyjmaTL3DN2Tg1ugQ97H/MyctccHxXp3zDfyHz/2wmNo7iNtlRsZWvDUBzE8H6p4S/9qmUC20jc/
j3yP3hDiH+Zp17/hWhnYPFMekHfwm5PvuknYrAHhg30j7x1S4s94agYgW9J5LYFsHVFMQuGDIQhL
XiOOcLx8uuorD8fZMLOi5X4JzuwFMrJE7XzkxNH6r8gOJ4CFdK1ELDxRYnNahqt3G6pBwiAjDO3V
jBDNFs6krg0EnQgOcMYLxuLfgeGy4LT9IKbPigLcq/XKSV6jB8F9X847U53eFECthJaURHC8POtZ
nOMUZ05OhzDQlkX341pVJh+tNXh+zCoG9fR6Y2AcNbwR7P/aKA/0Jiw6lkewTPQjowQ9QO9i2zzt
pRvzNsw/iFu7sfUuwxnRcuKT2vPTMUVZpHjIJzWYBLkNcSD03ekRaHzn2/eknMcHXX4s/ie3sSu4
tVevgGGZQkFgwn8f/Rlf5NVEEH1ij18TdM17jlEE0tFiJXS1qIvOjgBRFixoDcUBeW2/eDqEZep6
k1Pxt/JhA9Gyg3vGB8Xe/Pek/NixpakpxmbZBBwnfdo+dIR8nqi2mEPFg8IL+3Fsz7Xg9ULSgvBj
f7JdefaFweo4QKaav6iyr7BMpN9SGNHqaSRbmfdJar0jRjibWueoheC1oWky0Wn2NwmW4GAylC5g
n77J0ber+B4GlfSzxm7VNyjiA9RFHZNufekaui7WXNDSGhMbOfMMs4EcT5Zo1anqODbgkdI/H+Wl
ViQhg7eMevdArO7KW6cnSny4p1VLjwlODTkthef38hCg0RTEOK56wUIUzkp9iBX+V63c/zps3aXs
tUOyfp3xGLqA4GzOzHP/NXREeesTkrHABU6gdw3zm1Vo0o+PjtvaM1EcqArLed6dHrWX9WbwAdFk
zS9jh5IpqLxgVtmI/xfydxwBhpu8b2jbNmhknFtBSlX5geFZlDwDTsEvKovW6JXtPPYoaD6+o8OL
yeRIbwt9T61SqblHJj2JmKPf88O/u/ANH5qxpi6pzEGlm3uztJjBIgEMp9cEzeICI3HKUBRDuCO8
H3PV52PghyQfr2I6T75Cnhs5Hefx7bZdD7gUBarCpKu0UhZhq4HtEDoNCmnD5ax8J9w1uI6JB2gM
ESLllnMbl/RBtedZHtKLD1If0CE38Ici0LgE9lQqY499CkhyS9HGcUpru98niutM/NpjvySOn/nr
peNN0JCzTYzWqlha3s0k/qYr0I1occtkCucCAKLKcBVDlKbbFxGz/+vtWJogB6wSImpmHlQGpNhR
IlcCR24JURkucLzQ5ckDc5JBFG5L+wDCeWWDzl3Ubk0YqvCfPrIc3ii/EWBioSkh2i8AptQHc2LS
WtS3tMUHFThDHG9i4A8c0CmDE7ilxkpIojrqwXN4xZTiTvxeMi8IpgkFHtG0yWLIktAFypAoYqc6
6zc1aICC8kpqc7qSPP+c6ywUbmkw5WPM8/EbhTEQQ6iZSFp3MNzJbKFqu7nA1ZqCaj917dVLRRyD
rAdyU2YcJgliuLUWyvDFDTV1Y6U/l2w8+k/8nLotSe3WIJ7FZbXAD228+ZvHDv0jQ1VzYKdsW6vW
7r3NLD3vUKC9mDn6X9zhs616BXop36TvIOlOy4R/vzzleEwIy3XhV+t7zuw5/iC2tsxQtP+btAFN
BP076Fgj9F308OU85BXgze/4HH9+5Z0170n1FfAczXyiBbHk866jey3wS6aCgt+oJAKsYYzj9szh
mlffzsR3kRcgCheKPlY8G0si40POpBAOemDdMhD+Ej6qZyLxkUWJAk9uT3L+x3VGoEWAlf6E63IJ
hutcBnNHJ+5k5Gz3zDJf0KQFmYgo0b0DsmpJFn7pENeQYwpyMEw2wmBmwQtYAFpwevrdO6qHA4Hs
RTdJPiu/LInGgFu9G/CLQEMZYokKgY4T4HlsNLbwPDixAA7zJT3qeZIHJ/pODOVoz8dm+mDeawhX
njW2+XIs5kZPvMZi1w6ppKN3LiCeTPYn5v5QD4zwUn40Ltutv1hffZezfBXT2a6p4D6DnenD/Hyv
bC6HV+ObJOD6Fmx0P/bjmndbjlicYRMAeJwjrT9bGhBoGDcxCtqyurhyAq/saF5hC/+Dy1NewsHN
+RE4lUWkkEA1WkPNqbBHmFeQHF0JMLNdptnQbfP03gwgQyOP8mT0OgT0g4S68+N6GwfR1O4SDt9g
9czU82sbuyrDpRzHXiJupi6cA8Uo7DhQYAZhoOjVUzyzg82vFtbRwd3ALz5n1s6xCXmDiG9UXKZk
B3ukUDRASea2wM+Pw+WuVrwqxH5t1NJX8lPM4Fzc2kj8aZX9mHXoTkBN9GUXOn9LGZ9lHC4e3uS2
0fTH/DJmUy52hbUgxiqt4bXiM449XSwVrvRT6orU/1vDX2Q98MOLb6KIPhBwVvMim7ouVvAhajkB
zhtRnHNY5MGFSMojyXgaVoZe3/ofWvuzp0Ydrw+FoK4EuhvdIophqzRmbOaLKoh8EnknvAvNaNW3
gCy49uXiecoItfWYD006ArlAmuILni+yAPFGmzsw76evXBqgqZ6+eBTyabSc1dv5BCW+DpnggT13
SvcEGJJ2WlgfFyMLnOhPenMx+Oqr7WdH0Pp9R5mUjiJEpbmTT/DJvfsJExdVbs3OhjO+cBMIXZQ+
k/QlpSgBiSm5+s6XK7hq3MPP1EUK9+Q13/VUFcnp39BRtKAs8CT2+AfSViUTVXNSMd8I4HRfIWG9
0Mnsn+GX7PclmBm8s63LFFMCoBK8DBj9hg9UbzK9PWCL/GyL3ZElzPdYlGBoubWG8zlEbPfX11T4
4oMcY9ZgqRqbDaK926Dhz2C8jbEnyqoUqNYSc7zGBbr+Bcyg7Tyu0370IfxNb3Foo50K7X1rUEAj
TxP6x5zF+zQ/f9HkINq6oWLpPUQuBs8hEs5bm7cLsnb+5IjiVvoBxzSuCpOjvHuU8Ns6cyVLLa0m
jlFD6/uNCqKLFZkEYeRh5FQYZn9mstOakbgSghNiPS+CovIzuLy/j/WDJqqVVF2y5PWAPifKI7ub
FXkrGxpqDPOc8sASgp0rHFk+xZoEcwBJNddvrwSLX0fALkAP+AJIvUW+92DAdV7rolyQVHTwvcmA
BjnGtOVWqGUViEjSdRxDoc4K5S4sn9yBGvDPAvIWjaM4fgqkDko6/uYsCXKG1iMy4Xbm4SKjiQE1
llsOr12wS7w4KgeP8Al1bDS9AdoI/5dHSszs/v8iSS8SRndA2zBcyFB2x1/n33nx6ehPPT7ickAR
06cu8lIsNFCZWmRmF+/r8VgWyzh1hDK/Cvjp0JCHonXWA+967FxAVjNQsXxaGiUSZWbiqI/esJCb
aDiUB17Z+npOtsp0AIz2argfMFqrkJivsyLOcwHzStes05sL2pE+Bf09uH3wiPX0hLeJq+t76OpI
wMTOd7XD7I8es/3y1+WeIjCS8d/2GsaqkJgXKBlQ7QqR0skOAfywNbJOg4A0D0n+70pfbFSDekRl
yWM6pzMSX+S584HvNCRFbROk4J34KbecdEOfxT3Xy+TB1fd6/odflKtamRunbBNSOrAXrLHeb5zj
/sVSXzSts3wqN+2zvMP8e1f0jgsGrLUJwaPjMJ/WyzPipAWIsZpxuzrPM4G2UsxomPYUrqocLP0N
E/cBAFjCU4AK4f+mtwax00KPfSO25qANUJk3v/HDDF/GM2HyAeDWxap0Qex5f2GaBqAfrsmQPj/J
TtKji6lxsJHcqzDdOTKfMpZBgn6BVxWMNL3epSx7iBWMU0GHseny4SAeDdvzt+TCpErCN400p5F9
tXJineCGdxfkEIr2Nlfiw+t01WnbhILYyznGIFfUe+4a4O13DVWXAZQKjrzQRKDfk1XxQQjL6xEd
+TZNkVTO4YJyDajtqzwsViChkWuDCLygDbikBibUxgrEInVtaERrIKSPF2wi37eGYh8k6xJhFQhD
Z8av2LKF27yvoWNiGk7O1RVr6H/k67mh1+kH/NupEkN8s4FUuzLtHU+vTENLEn7A5jDDMqh1YPfR
fWHPM32evimoX0WAwZni6eFgV/QlokOntF1enNFbJRp2RSbVBN6VjsPJzR1VlGNS5jrFyjqnWIR/
gdiP8iJY9tzem3kIJA28EgW9GOfnKyKoHS0PYnA1zgTPybTL8gQw4uiPVZ2IpbAmIv8i9KbJ1Xn8
BvclenenJAx43gzQSkcJ994B2GjXqbWQotdLeFb0roSzHpLr8KUjgTfZh+GQ9dSnmNwJQhDLDpc6
VwtZUjniRhjTkbh+iYBqJWrJsmm69doFY3NnYKlsxxpVmi8dOyb6ho9THzKeeu43E4ockg1CZ0WP
0sas9iNCLuVCJe+GloP96k5+tmzfBVDmv3/j+M48+QUADN3zl98i+ETSPKfDhPGP/uTJAVKiIVGL
uHjq0XylB+s8dHrNDcAj8ArKM0bj8WmlN9r6JcaLgWKhSnfgJLnK0oDuhWtHMsNIayWsn//tYItX
QKApUjGWrHWbC/y944qbFvSTDd1q0B9XoZzdh/KYjF/xubj0qQTuwDWXuH87Lgf7Om386GyGMfw2
9fK/q8YgkRWT+VtzkLmAegD7dHkHjrIvk97wtNXeRxohSAGq/65F84XJqliFa00sbjPXpT/vX9cH
o3G1TZVX2cG3dN4VwpsAjEm5QRG0TukLhyG1tIAc1yXv1yY6IcfLDJJW9pVlWMEC3yZUF0VVEvRr
gohFlxa9Z+G5XEGKSeA/5q0Z118BSdDQMPtZktJZYcglIyV1ptK37Llw0hBNVToVG+EgcdsN5mxm
s+KizFZnZKqvIZSWlgN6iAWd23otaYuFOHIbui4xJ+TqAsA4ZJIz9f5kk4BGP1wEfpifMsNjwX6F
S1SdlBiGPFNMtL9jQpGae7TIVj6IuiL2jxtvTtHM7VBu4TiXxP+Rmv+4wUzR3LzfO7jGmmMEYM9h
l6vQO/DphkHgNb1BYeHpCUHJuLV7TLLTHIk7zKKP8tKVX9OspArfzaglwY1YUjWa4pSup03uMxQE
dUk33rmoTqhqsQ70R7fiaeCorrH/aCXgwjsfJRmXAjLZfs4IW7NvLieTtWi477WYhBicoLrCFr1U
gmJvAeXcK4MxKAYR0Tv09UG14pWcZavHdj805dSEIzCNW0JHs7fW+qNJ2ZAg7aoXQJY1GLqGcIAd
TEk2oXnxdCiJBCMFEG3KV/ffE+8TebhTbfZ19YN9dvB31OO/nR4rXn9uRrIPkbI/cVTcSMxq+GYi
rsiXeYkvixw+V929MwAF+bflU4noAbF5DfAE9Y1aPWUk227BsorcfkpcBfLYoS86rc//PnQiWbyT
TT8cmWkb8+4m5Ez+o1NTJQMaCbSLsWAZhTs9G8gkfAbel3M4kkAjgDyTpJxfra1KY9k0qmXl3Xj2
rqETFkSxER/P23cUk+grPzRkdaOwWwbUsvS+0hG2CG3xDrHweWmccVXVxPxRFWOFvV+xn5ifA1WG
XghTdWfAi/ZFFzZUnJNuIqh+4Fe4NGk1PGjIR+zTWqA1uHhn/H2XzRE7UzfgsauVIaof3E6L/mPP
Peui7wfAcgZ3DXl+fdLuYziv487uQAsa0igzBOK3kP26HHb4EgA03Abuwgk/K76CUyS9B3esW+jK
GpaVFYSjSEVjptLGAoFJKkg2mcyoKUN5JrF/0EXKJWPVKXs9FQjTww9aEred6gCAip/WQxyz3A/s
RQBocxvQ+Bx9mGLDba/u8vw5LSweSdkQOM5re/TAmzg9HxFlo8UCxV4f1/mx/fGrkrgs/VCN/Hu1
8MwUnSRGMj6CEUl7Mj1c2WlarJKJwcgSm9W0Yzlgsg2CFKnJigSgsSUKFrxWy1m3wOZaj3MmuR+i
7U8aIX+asc6o1mo4DkJb2tlIB+S0XF2aL1GrMJcupQJZVOoEKC7SjIMEF2TcZ0TpAiUHcXXVQYjf
/rdt2wj/QlW75pJGuUO5+Tu794Sh4ZX3pGi9aGDt/sdgybbmm9GCgIfIsLvGOQyjqBbleYZWj/ce
wxfRLcR/bUS60qVX9VFYBbQN1RYrzLojnBae8nWRsGHhdj6Tcnr94ZDYi+oua3TNgN7zH3VJ3FYN
jcWOWc5ytimnxUkxWhSXs4gO37mVWTYN5FY2ZUIcgooeCLBxxQf8HZr2Rt+5RWSTkEzvt33q2+l3
clSybyv7CwGDSMiyZisN7r+dQkb58+Vj3soohEZceh0/ZsZfAB6ev/K9JavrXtk0DyFDtDbaKnu3
Rg5ZHryX6sStpcs4xvaWn3d2H05rYulRrXBdKrTULRAgk9pl1tEDEweJYEo+Cnu0WHyY7Jv6FzzA
Snk4XwwrIRAkqmLt4Kf1nwIUjM/SzAqTr64YaGglWH86+Wn50MXHrjuSWycQElj/HAG9a5GOt1ot
hbcrw0XS+k+mUvOl8gtciI4VIHcu9HXbdwLXvEp90FYbOxxK6MkoEMoqi9r7uPWklYeSg9yLK79Q
N4+ebYE6R4X/owiVPcd+NVhG6Mih5NI4jNIpwayjp+LkPNYVY1jVidcldOw3Pr1YfWfBY6NNgTRH
0cmgUW6miIQ1FbcxMjN7Mn3MGjWwL0Z/rsL3k2dr6jYuTBpk28jwqEWLnGdY9Vpuxz5TtTPal0tO
SB17Rqhp8qXnoTgJBSVUGSszqMjnz0a0ZEBw8BMkUEEL34LilXSzc3cYjkLwYlrgulKn5C8Mmbpf
mvOHUVFmKy3vGdfWi+sRWU6ElDS1UHoy2nEL/A0aFdfuXNSZs51obwbBXnL/j+PnoQhIzPnAfHo7
iyddzU4iu8HnHlxatWE4VeuHzCSGVgfFzlHrWi443C4Bltv/rKOp6pCHblDlMcOwwniWh333mY0L
ejL1pq/LAoNgsswTMt1NLjlbIeRVCZi4cjqWXbCLHqfGEZdkcSwNTHnAUc1eM1aKwwo2EhAq7rZ5
Uek2TOJp97kI+T9apxyxAqq+7Vq4KKfcrGqyys+mvckziTo7+EWvRYpkxr/+HtEcij9uT97WWcmo
LnD2hGRg1UOYSMyhhBQ3UihesJnyvP6DLs6BCBfzVb+CGR++j5PB+O4sA/H11ycRup909G1LRnrf
Nd1RKGwT4PIxuaDKkl3uTzRao77p/yZ+KujC38CQszknQyMETiTXyT6NOaTDVN80e/pRA4P9b8go
dlH6aN76Tkhdq26ygjGJYLcjqqsljBx56mhAWMyAlmuG8KeccyabsTc5cXOLGtMBWNjjS4ZFk+kP
v7GyJI2A/b5iFp8pmEHuPAcObVDeT9vJC5MpzRx7gH54BjzflbeEYPd7iNLr0XIYO1at7FFjEChq
GdQ+IbPvomOzjP4L+vbqwjL4M0d7qn6QNmuTF6YZnUYqJE69FIgMBO3FvIu8HfmHrQGP8ixmSoSP
4s/8/FzmTwAYcSzWgnpkOURL3FR2LzYOdOJI27G6aUCWoGPPzu3BxnEV0cOqVIdTg+XnrBKhvSPu
y7IAHtQALWrLXzfUC57StS1/j3Cp+gYOrkhEwA4xFolVlUWaCehsTbB8nBGqHPAkU5LdhDrA9ft+
Bc0GTOoDpetG5dvS+nqbP5AN1tUn5AEXPPtWMUmvnOCuk4XA8VL0tPKajoJh+uxu/Y8rsZe6e62Y
sd2GwaC4mJ4TpoUOr8I3exUB6llSSnT+7B+lc318czy1FXyvpsI0ulEOIV+et/aRLrt0zQ2Jafrx
KapLGLjK9SD7+iEIp+TrHQ8XD4VoOHLey8iCMv7EhwnK6vi6ti4/Kv+RfA8VEeUSSTF8Dd7qbWdZ
nfH/EeyvWVfpxmqiKexqq+ZDDp5MUafQ1l4mJMOcqX9/07kVcRMjkmhHdvVxU70amJwqLpR8+5+g
t7ZZ5RsWNWiaMoNMqTTxPIQrfATTIc0AMN5sf58JZatJU7cexW/LoVO+0PNWUgPNgHBV5iDbg9EQ
wkNGD/HKpIVh6afl2Nv8VQLFLdSR+kUTqQ2DhhK13RQAZPHuXmqPQOiWlVUegR9JDJyiERaZOAXO
Pxhtc13hhIKGv0qJjBOE4BBhsJo1kNAvmpkKF0nNxT6U9l6Q8H8TEJyOYrqY2PexeQXYr6ejHFFY
eSsdg4Tl5+ACkJd9hBUzROjlep9c8ld0NYWnNloZW5G/hrg58kJigCDCpTnNitIFTnLX4vKwp4XV
DQLS3aJQyib7GWiF/9LxoEE7JLUlMF2JIGAb4kRcffHbtKST32+ssfQkGLPK0pVAl75K4Ly9sdwH
uhYZabfyIPxcNlay1FZOrwllUmDZcFwoQzBaYNySjk7/JdCTO7PMZpRXKAZZGCha+/YAJWFnfERA
bHHcG275p9xhqyZC39Od8NGvtctMQcJGNHEJXFyDhQv1/niFrYpApQ+O0SfZnXuxw5tiJov+KFGR
oUsA1MbgAwq8wyx6y5sFNYAiDZkE79s9PXuAhq8zp3nQGgBxPYW3cb8iKo15Y9m1We/pAf/yrYR5
RTt5A9Yz1Z6q0oksR4iAgYIL+TnHD99rjFEGhsuuRwfJTz2uNYXQWqTxRlcYhpQWKE+FJmIUQc6i
Yiu15JcDQfoAxymx8Nb5a0uD/C9kERxv6l0ULzMSsV56kV7wTKFeHdhpWVY6cdRww0fwFl23rHQa
dr8xsP4T7Mo3kejOUWnHM1Zp+Pt+MnqJrh2947JFHv5+AzqcbZHTRGuIhoqBdztydEGV3AEiGl2M
fH/9OLFjlZyB6oAL9mrJjMvt4PbGPWb8PYzyIxc+evKj4IdKjAO3T+7jt4i8WB9SL/dVWI+PrbZs
Mcxkeu+Hw6wSHcsZ3s6c8VGuoWgYD/gdPSiUSJ9V2saho3K4Fn4tXogo5hueHQ7LESArfHRvHM2A
3hi4H46EJowo/NJLZQR0k6/v9RK1X83PoopmvWrTT6d0FCwwgTeYZKpLDMhZdNvL4n1Q8DClLoI+
yYGa07uIpQbJIzW4TrXp2UqUdb2SYcIzaaBPMzqK+gUDVfmgt1n8PExbtHnQnEjwOJGOpEt+erMQ
47Erty/rgaCUfAs8lxlv4JnILBg8vFxrGK0aR5g/24GjcGDRs9RnWtVcprPyofbiJqs6e9mMRpP3
j4o7QDxpFEREHRZXp+iwUY3I+3M00l3FyOBTWfTm4h/2Ab2/cfVqlOqC9lCoCcff6mOcawG6N/6I
LBnND7jFqV2dYL8TNUVLtVCj4LU0tf+x3XqLv3zGEW82NnuBhUyqyW2BdlkvlUevHbe4oulJQcE1
uNhHwm2iyRxJjcAU2kH/0htnz8x2LhzfQFEAPz6zRsQKzIG7g3VFQneMMj3iPIKUbX/ctjBCkBhv
/lDrThEGWD11WKNhJDaxDjcE+o7Sw1co7CY/AexCiI9Vj1AtKEzJ2MEikVq52yTJe2SN/g9Q4/Sg
5xkO2/TYNuW0Mv3zbUzvkBw7w8jKZT3wHWoBXOQzQ1Vf7yTFuMdFoQmnWejTvEqVMSCrRJSOwD8g
XIauD2DRtzVWw1oj+tlsI4otlraC8yTz86q04qEum8o/ga6O8WMmygPa+XmECRUoy5uqe4Y0bwvh
M9QuCfiraOwhjpcuNN077j4LL4CsYX/lnBjrVZ9ss375eyHQ+7NdJEXG4rNx683fCdxtI+kD9SXl
ZUrrXiNIQjXzu3kZM9LtmopJ1kzaKfiXX8HVx8MiEIxVvU0T2Ku7u7nwV6mF7EQcgVTr+5n8EYBY
q2QZqu9LAYLpY99LZhVB60KSSzRAGO1WUf2IyTQWfkv+x0zViO3I3NjBpFhPcqe53N7D7WNjccKx
wdf35FWZGFCoX5Vl77bHyOQxz9DWr74h5pN/6li+tgMNiMa1v0lbn10jzHpL8F81r7GJBNJT/8aH
Y98f5sGh126qS7O+ZLgCZPbrtAQI9UXtx+vmUVTzMPBg6sEsy1LoiSaDDDzyIKBhsTxR/u66kgVl
AP9MGbbhJ8QOGQZvSGQjDuiytavLJXdCr/LbF/+wsxiwflmYnJ0ztba3IykJvfIafX1OVbZk/tYH
07wWbX6kKuHy83fCLYEqbTfUyKTIu1dhj3jyWNsEgGTIiklHorTibdqBEw3DmwxNfUOz5pzvL6+f
O5DoDBI5Z5QeKHJhNqyuan4AZ0XrIKJUYYUxbMcKOvtolyfVVwPIU6nUCci5rllTgJAi+fwh9IiZ
Ih5mvsC/nHbZn37TmkJl1k7fDyqjw4PJyOWkP6/A4peTEsmOfRycjTAHqTj8uDx247qli5PoG86p
pFjl/oZMmpxHIgz81gbHwFykMx08nsTOTXULNkqgFrQguopHYotU498lFegCUWg6lALoPcKH5iu1
GqdfZs777pVVoTUQ/raaxIsRQcO/FbRN4DB+YjyvTsXeGy8V7OhO8kOyzq3cm3a2EgIiA9LPEShz
VdbRueqchJFHzPZv9HDkD7T63Q3ZgVVwjsUP/eAsOHV7f9DDmH6CyKvErSMOOMmTs0uyUiv+KF//
pCf7RbGY9/a4EUkFv+kPEPDDoO4g9EVue8lV2NVmG1NZ0v9U7lCddSM3t689+Zue3yrXw1moMepu
ifBVN4rIGYHrhg4beYTYltQr4KBVjP28O/qhk4lGV71gwPSj0RzbA6awsCn3xfnbg5mOiNaDlniE
UZ8ojzTYnic3PCJxRVYCTVV+31pqZlY9ypET/9q1PpdyGtUY6binEfLNtp4+Gc87W8n34k7UbODJ
R6nT12/+TGGfLwD3NBPiOBqaIxwYE9ZAQnhCFjgbaSV8oGKqRQOhJCwmA7vWYFdnG2q9uitWcAor
bglQIMapWRx0H7wV7UdUjbYqGhdMaYXRcbHErqr8swDik18yAYjQ5VMn5AxnPQRsQrwIV1Labviv
dxARhnL96wLcAgD5iDz/eyZRqQ397XU0uxwbk9oRBeXb+yiBsZonWG370GMcd/5as3h7uXwOYmfn
bMAvcEhaA2KDrhBURbuB0tlBtYkCbHxqr0X4bin9k+IWbiFe9FtUu3sEdFeM3+ZEdx0vVdm7Ypp0
1OQYjaPbkWul7IetOomuMgORry1A8OJ1yMJFO3IanbFMTnou8lr1+OccskPYHrvqc/3R8seWgwf3
5+VgHSFg8ooUHbK///9X89BHAygmjbVw5TxIl/T+d4ytl7NhNYcHn93YLoA3qEmFuLkOCDgAbhxw
FkHYV8tyyNl4ud/KVTptPvbiRFF2kRtGCtC4XTtzvGx77fXjM+FajZmsIPYovXVd1QtTIdrK2Qbq
BXG0KPk7kIYmsP33brZ7/4bZLcB8nE3hquH6JQ4qElEDNkhZFyUW8rFLHoCPn6cioxoW7wA9SOPT
61eM/SDBCNl5RH/+fLRfFLXgngMzUn5x3Db+ehMm5PJow1ekf4iFcKjGEwpqQD4uUwQ4uqg8qqvH
saSXyMrwXmiRNxmF7wWsuIA0OCWWRINKObo/OI1nyiPX18VXyc6mVBe5w3Cq/3mhqgx1y6Rrg5y+
NQ2cOpt9CbGlXVZuF1os8gGugGniReiW+54XOmPsCoG39p5TeRn3oy4YlSSKwrCfKMSc2OuwUqrF
6xKUI6ix/+No2ZmDVhOuBCZi3IFZFSvTyABf3P/g4ddQwxhlIbl+Yk0mv7R4GE9s2gIh+iomW22U
Qt2MTmdTLG6i8TbEXjz+E0SHHI9KnOazDQKpuI9AleEzDHtmL0HBct2iEdh43NhIAOnOfZIj7UMX
Z51Jw2aOc9Mk+ntHmGAeF3qW+5pTe2IPL21ERn/glM2LiKEFXaB09/1VyVqnIXFa4ksI1ZdzVLdX
DKlEVECl64InWvw/rTbDK3sq+IgaWZIXoIQpDq1g0IljVNJxOfBGU8/EV1dvJXaq2SAxOsJZDOR4
G86pVy4rjAH3zZWWdx3120MvOYWJulHuU79kuGhqjOlTLXw2xu562eDxHx8uitlRZmTy4NTJFdwC
u2W3/cvNIRDAEQUlQQw4NStfMe0L5/hHIoUud+Qmw8KI9ubNU+VdqtZnztKeN2h+xc2BsjhyT+1c
cGHppzAFEYRG2ryZ3fppoBKOcmLbLFqZ7FhRmKT6A0FUDwcuFb166ffbp0UvJ7y/nQCIWxbR5ep0
ukwlS3bKhc5q2lVoPXp/nNMx/mMI34Jcp+o7XdXW1pjSeOz4/2zweFyMKW+oGMNgCHAtUVTZ4eBd
F6QWF9/75cRrii/HVMOQGAxyzWsatKnVhXePcSfxu+ZOf9od/+KGGbF2Uhn3nGKTC0C1vkW5faBP
48a0rMqWosy60gLYUl2akqm+9E4Z1TTwuPreQhThWAm/5q+miALcCGURCr4MBESUPCTcYMknbkPN
8Yfhf0U6cK+2gKlKujp7fddP9b7AtVzozD+141YC4ni0aepxbfUO5AxPrHx8kq17RF4SJHvfyY7a
bbIKD0Uy6AB5jjSTSdoygLtY1GxE1B2FoiJXTERMF9yHBja0iqp9ceNnnQFvPJfKNJ9378g6OFeV
xaIhZy9ZgPtHv3MluNIGfOK4q+UZO9wdlvmLpqcjkM1x2ramqux9+TqrHYr19SFihYFIdM3UkAkl
N4cuuQn789PdY320eAyvA8O9vyMz6kASHA8ZvU4bJGyE73QEJrPFINVhaIz8mv932RSGzO/ybQVf
icW4nAtMmBJyl0lb/nZawdTwzzVH+5SuAXeGwN22Ikj+GEaI8dBmeR1B+CJc/g/tQFvvipgNAat1
HTNTRwlFxKN6RSQPHswmQ3B6njwDZQd9ZqEuuPOX1rOQTr3WNfmVurM3BeAoAJbEZicrt0Yqdpam
ZaUqMP1t21hv0FTafi32XvOJg8EhKsYjXFdBwOjOBJ4HiscUZH2LRM81fRnZ4velSpFz5A6TvLOB
nsjX/bn6KZ9xCWMfh7U5E1HeoYrcbQKTMP4xe61MaTxF9XwNlxP3afeYk4zwS+uGuFkkqSTM0zWm
nK3kytl30DNQXAxKpL1SvmGZDxK1///n05OiUS/G4Otffoj3nBGcjGAC80b4lhf9WDEhwjNpTq+w
4w1IhAFy+73FjEG1THr063VzO60xqbnuewpzLIy1ql0PE/SiY6xDwd3myIarejgUw1/BvnnpYb/6
RrQgP23EvAtKGTGapQ0AdjYp1lQcAz9TLhGCJMKJXfCj33sbfhLH58Vd8MwSD22SQmi3SvULaGTg
jq/9txLgn/PEVkRxZotUlsxmQyjcakqgzx9U31hfSxiblKnzi3diNiVQYIIMOkrXHjEDGP+q9ZZJ
9AJwajjNb6ajhqX/tOglbTwNw+OYpBvUzNQu4nbUw0avV8fzJocyGeyPC/77m56ksuDhfA9bLBPZ
pIs6w8E7oPsts7L0ctwlZ+2eKPwfCF1vXSofzfmi2Zlke2y7fC+FmQNus80hSZ3TYB3Chy0GXgDb
OhGmU0H5U1RdTE7Nqi1FJgGyAJZNRWXT+cHqK9Q6RmEf4Hn4HxfwACReiGIMoCnVJNeJNzRrDj5J
rWrz16s6gCk3g+Usm5+ftO+o3I4qsrRw9H3UnORe6/UZmImov6u/Tn6/boQhJPlW10HKP7kxpNxv
8SzItCVPi31zvItd4xcWB1KuCuqIcPPVcfRShYjHGqB+xDkcj289UbQOK/JTujFZmDt0h+W5Izbl
fu3RCtGKJg3fQmp9c2YYUOi+jbhoZERiPmPlkRIreLjRhDTwwM8FXp57PGEyqicJAXM9/cCOvYb8
hNUUk60dLAha8atoz3u6hnRAne1O6/ilhKPvN1pGso6lBE6cXry6QzdiAPs1cMMeDTovnQQT1Ftn
mu88N9HNvECWkNFcHbVMiOpHl0qLGMIk+kS97H65ZlQ5pfld2MnGnAUPCetN5NLytuAT2QZichPy
SVQg6s6zQkfTHzijoKSKhVga+0Vj9YtPPOOteAcAT1ASyLyQx/IMv4ZhKsOSmu7//MhiUWvQf4Pv
AaTzb0DN+lIjz1KGEqMl96XdQwovwbYtQkfEtTZZf6yWoqzrKfS9cGjVrST+PPJ0tnYSyBt8OL4I
OJUdj1iN+cqJxmJMH7VBxGPslKTvqb1rCLx05xfEcv1IOMkJ6XrnHP2SI4AR0fr7PY42On+hwqWs
9Ai+ZPRZqL+i3mpGr/t+Z+GRQpqVsk6tWHk3REJ2RmTa8rEuNIVdjUapDdsQiD18wSbhBqkYXzN8
nawUJ+nVrnfrFabHyA0CudjtZ3I6oBQQGDdo7hH4BC5s7uY9fBMs14d2QeCX78s2PTvZx3I2ZVIo
VNbUGRjO2wLbiQJE2fGtbJ0HvFOZfOxtcvMfASdsMVpX74JJWnzJYEzrSCOgbGYzPEv7g8vjlZq4
QsW0LNsWhXo/8VFhY/Amw27wqwtspigMfsT+4iHdWDV5ouNIOJxP0H2nDg2kLO2zb6aWWB1YS1/O
qYNW3FnVDvuN55mhZk3xXtSRAYHv8IoNP7vDXonFB1xSA9uU03v1FP5A1uq0qByBVaglAY1SrLDY
YqO0Rwgtvgvp6e2oWjhXl3SKRER2kF0I7FzK52HO07yzzyY9MOp2hP10LW4C1GCwdp9mi1AXFsaD
gl8RlEgbK6uMALqJKII1+UrXR+3+qGO/gPLUhH+A3FxcmiqJ9c8k2aoTRqp3yaMioh8B9pexxLwg
EoYFOARgxUh9VEjr9nRZ1ooHANl5vojqemUnPKLhOJpGbZlT47Z7SohClFw5xkPsXSb5m25xuF3A
PjEEgpN+vKsEy20RQ/ruaqUsWielGSQq5hMle1vdyTneQGFCl3INKsmDFvKgPa6O3MiEcBrtAPpQ
xuquZQpawbaW0likGOtGWJcrI0u7VFL4KJbS10iTfOn/yNLqAtn88zWRRsvcdlMqWMSvPr+LSKnP
BxJOp3VXEAw+EzGgeSQcyndEJYioR86ZaJrsmIAv47qKQ6/cEbZ8Mb7WbRQGwMU/PttIRS+0IuPX
4/8CWfWnw0i8h54McMKJ7X6KTgCD58zb02nLooYxTi0g34kJrfKvEq6vdn/YNH2gvLzhgNbwSCn4
OLaXau2P1ZM5ZLvwX3Euj5sjuwgJNlaO+13mNExJrxTT164yROFcfnmkt1PsjonpSqduPwC3HM/W
FnXq6S3bDiNarWpSQwc8JV6mkgHIRnAK7CshGkQZNFxep8WKGO4OuBTHGHvPPbgIejPHdgY5V7QR
Y8JHQA64wH65HHVpvkvcAr2GfphJ8qXbclYDqKdfIZJMVlDFrDRaAEw1ai7EE5YYLHL2uu2l9nri
LgZbmhSsoQhK0DfjAvdmxti8ATD5E3O9jFpBPSKOwYwOM/oqYwESpHoubf3OxIRhAyJ6IaOYOdWK
dDE95BUsWO5gDsHtOEhKdvnU6yJknn+iWOPftqXQTzUZlcnWqFlPDRGO6DArlx0XSqBNxKDZkvhi
n+LV0TtqyuACGYVuuojWvA1Q1RwSldacHdjKXIqmPWvUNz86nftEgpWQghhEXXuIwNblo/AkYgYe
aF0NuyzmkngKyGAGwi2vrrE8dQ/zIxWl80ULPfrfYD4J6MSAmJGkcPyGz7dY4B+muMZUevwMuooE
sJNjZM9J0UyFG8mv6s+/UvSTNUFjtfz73UxgP88Nu3leY59OMTkz50Mf2R7EP8a6YmsFxNc5BuAs
SkkYNUbJp4CKHZDW/HuOACFunp8JFvIFNC0EIiSHv2aBhoc6FEGj0TAEozlWfMpTeAXwTNgwqgr9
X89s19YXSgEn0ThcYaRD13BVf+Avlm8gml/qVhRN0wMSa9Mz0VmGCLvEcZU7DUwlvrtIlQPfwdtx
+ngLMXmhIhJTe4oraXiqKgUj+NPG507YpIMTYMb2pkedkeGzlzisjomnf3WMGrn8t0QuGLXyVPhX
mnMuhjw7slg+aN5/lIkfhV+e6WjKwW8zSk9wX7hikBzeyKyd1RBMmH7nJd7nbgx8HTK88bNT9JeD
2sQhGKGGcTujSiwfznhyn51BPd1kFOxBYbrc/FFsf9PeME3OfoySU5IOEGMxgzWcYdBuP/y9t+G3
YLxnS7EV0E7zOr5yZLAoYGHoqkiHeKRBbY7RVKQM5ZoUHMPj4dNkYB4JJv8iKnJPegUfbLEKPCRx
5xFZh2+rrRXC9zAwbk9uS1aP+r/9hztuKwTzT6YqexttG26/s8es61VEdRjC8oT3eYdi/lYYWDuL
x2myi95VF5tsiPddxAGm9m7u8jkab8DmnUF7D2nt5Le5gLAiY7VCLA+Wv8Cq2D8zQIsEik6B5t+A
/06YsFoRdi+MQ0G6NroQbYYhdbNfUvEz8oWsRoK5fLpPW1lbntexNDAOgPrlIfH3D1uycbL1DE0e
qamLYgCNrOHalM5kmxp6kBayGpJwO2HGZHewqizxCUdoNYo3l+8PEd8B+4+uwqDDYnBh1VMrCoX5
DLMc8kuZXdibdDitd76g41vbEVSenMdcmxlPDt6AR6pi6HruyFa4Y8kISJSGw1fh4WD3u0Ru5+e0
KCaXtq4mRZtdyahbCiDR0ZfjZJstd1uAflwGuwTADa+744XeBjDzFnzW/Lru6myiOXnbZmUnO/0/
+mAvwtkXLSykJuFpfY6slMwGXqiIThkXs1hI0ATvOqZEFV6J9nI0feZ0lmbH7KpOFcNXVWZKB6ui
A0r1LjtCw2rZOtuknVFhr71z9Vtm1AbgpOZUYVeHTs68psfCZ2Uaj8XewIkTpT4wIVEvbLYJcRom
jgOnj+fef2JkWvDPKT5RnDlmze61YNWtY/QeUOmXpjD7asBXe5JfOcETDLdz5RFqBr3+7Jsdc4yx
0/bDjg/13PSIlFHpUsS0Fo/IP9l1sqgihZSCcxLo44FC1rx72IKqbd+2/lwiIw+K1qsTAw2MnnCN
cWGQksQS5vvhOhPPazvNnCcMZSfrAK/OPf9OQbYaPDjCJtIY1IP/o9KggsAl9DK4VxvlS3B0J4vz
SnErFW0rieb1P1vWXqKc+UqhdpJP+gqRdwOsrhQaM4814x83UCEvDFSicEXXE2ve+S+WOWGGZPm+
AhRt/NuZ6qR/R/F0OvUfCfYh0Yplbrs7BsUIyBn6tAquiWfrVL96mdMI8c+bTh4Dr/ZIBmmcl0hv
Jx5wk15wA/XqU1tE88+hNCEsj4FoLqKQY+gb/24JaYyqb3ir6vSoMjY6IPis4R8I17bm/Ag6MDI0
g8fAMoODo15aBs7qsDDQzheO/DTnBpU08yb2+XX+lEOzeGM+jIfM2r+YV455KIakr7XsQi4sGzEO
X4+YbeRQ6lSaZCgUR42mJF92DOc7/3bMI+MFVOCXfzBC3r0DzmY7q/xBzjc2zwJ80rFfZsFrJpS8
WGHofYqKWt7Wx/ct9jnQ2vKzGdJK8lOJXAkK/gpR0izayLdiMsCK9vhNiBPJdNBFac9cMv+FvguD
Jg00Wkr9n2IKNLufKjDQN+1LxQ/JABc7+IbXi6636RYgD0gM4eN6ErqKXwCdH2w+tz7WR0+1a7r8
5oMEni4N0WoEZHpfG/YPhS25Di6xtUydbMIlHGt8meM7QSXZlYree5leUBqvH3GoSq4ad0yglZ4h
y7fYvkq8essb3OnCqBLSnHQaZkACMMEu9w8j5gu5DsuSMAIBeeF7yXIo3WAYQltpfUaPSMhtkko7
oyp8d68zHigmupDr0VUq6/3rTthvR4tmED4Q2vTrWRvg/+P62TjiUU3YbnJ5WvjeBPrRdw+TXVNi
GuXd7I2h4iUgBXuE3j8tOrI9+19sQcbMNoctH7bfEucs9S1r/awuejuJ86dMAoTL0zJJCt/LuSbg
2IaMRbnVd2GxCjcLsYdPdS4IBEjNUeC1zPTMIPmIIUIjhEBU/rUW/1tHvx+NlOKmfwujWbXbzJEb
BDP72ueu/ioKgrzFKmZyYGO//QK3TtEGF2J3+mZvggeC72OOAhRUkq+GnAHeEE9/A5ZpCW/YRLpp
URw8dqI4U7kG30C3TCSgk3FPoaDRSK5B9EpwC8JUMUXn4UXfZMlnUwDUBlbCE4WZJ6oACXfY4PQZ
0vbkHbiGCW1lN/FGJ7EYMgTK/VT/uOr3IAD0QSQ4nRN9UVZuPJQ9FbzYGHgvZHb8c7Ij2SyEEOdx
CAyANtNCLoEPHHCpbJWlnZ0KJApCKOczeHdRENxPWh5nfFHL16JjyV3Ja4jxT1tMybI2WGH51IJX
VSGYnt6pDWb6bRUn6DX3ayOKb9EzVzwS789exmWcETqg1z3qkw2YpLhX4ARHihaVonXyOgavhpFj
WgXlY3DaPBpVRgJM+fVV+uK+tPC56GQhnQwUouV9YSO5UYHuntCEpMsaRExDWlf2TDFfKOjjEDa8
3bDLhWJgwnIW0ltMENkTigbkZ2RBJgfJ5j78dqNQDxRi5GSV4dA/9AtJ5AZvdf4nP3fSAgecoU4k
tQoocstL2m55NxvQ2m88Pbs93guwnH+qi89/XB3cRFxwdhdG8HodjAejhjfujCFIwt0uaI3R5IB1
E2+XJ8suFfv2nyCimVGwSeAvxqPKOfs8sITGctB3Kga7TJk/XNu/WTEOjv7uYTH4SgVHj88JDf2p
rW7jul/AIuGwSykR92x+Psd7SOWoBjQGvzt0QYBa1//c1Rb0sx88jOakoX/i+TkgOiAdmNvtct0K
cQqSglDghPN2sIVRcyJurETKv7gtNHOvoR0hJIhopFQyHrWzQHkzqU1FN2cSeaBsijJAfE3BnoZE
iL0igyOkW1Syzkk6kwASaRz9UgSOUuLI0kuO6DxF+L/swuZ0bf53Y3heYkumOdQOM1Xki6KuZ9eh
iRndHnYiML2aAgk4Qj+ga4V/T1U81Slnrus4IRKsMMuQbZvY39At+ozYvAU1wyBSjxe15tycJ6oy
aBLFdSF4ZMYzBk09/BnmzojJiKYb0rUjZwtnkeGXw4QEtrJiexh3O+IUX57W/8lcAHZ0+D+SLLvs
D0NxnIS4PRbTgVyX+orZkTrYXMVlbvVCCKdmr8jBKbhPQXF0gi88y7qyWDGfmb5kRxrwIcQdp+ba
0/xZanNRVtLdEC3GNQ+I3Glkt1UX27WauSaun16tYBH8QVvXzhXgTZhQKZo/vTlHX3aw+PVO6e1S
o1CODzMbb4pahBWxXgiTqGu5hJI7hNGznftHNnznxXvK+XbTHnoU4hKxeqO97dZxz9yVk4VTLfLy
t4juHWd+Uu4zwTG65j9PqBeGAK6RWs/3sK2CwBTcmzbbzNRyKk5Jr4CTsOJvkuqqeIzWQJa7RqiN
88DHyrgRpfjK8XYTnrhJMyuIuFwug6PC14F8epZdDyxGgPMQ6majgS9yn6fLkwCttEzCpwnTIhxI
BPC7d5wT71TUBLWHH+/iCOHymLWPKhzoOPBEfMYlx3y4l+YVeqwoJlugSZfL4XGk8q7O8bEeGHA6
/0ZJuaZmpZKNclh+jL/ahW1CtWAk6AgXv2l5GqqUSGIp0RUz7MZi2mrJUczuzcCzxXVQkcozmQ/2
AOsWohbMQybF5ADGm7oJG6IbwV+9NMKptc1TP7G41v3ITM/diP1f8f0drr1YH8LPVnjp99GkD7TJ
pPFmerzlyOA5+Pcsp0JHuCBI2Eo0uOqgHoYVmk6b6O0p6pEyw2C4EHAanVuATRGkKkvSVAp+daUF
E/9BWmj/MEBy6DTHl7+VQHu4A15Ec27pMdO4BOj6YgtqgXkHE6wk5mBFB3PZJ962IqRHq/1B1thS
a1iABu+H6/HQyvYZs9XjyEvKV2j/AuUwFGblrY/588V9hZx9DCp+aPq0l0Qi4f2legCxFTXI7fE9
47KQIkalOWzGP4LAwDsN65VzcqhOA5RRtYc7zcuAWTKhmA7ss2LOzkXcj2hN1cuDjE4uDMftFFNu
Q694oszgocYZiY77eOraCDepxTV6/R3kZut4TbA7gWbqrFEgqB146VVFhca643Q6zZZ5ZHfUdnEY
JJH+WUvjTjlMiHyBHhDNUR3oJGBbHobjJ89XubxfEb37scnNL5ni3GqRke0a4ofV0Coa219SU0SH
AUejsRPG67SLBggcrMkUCfOb4y1fTnxsvzYOTZvYKhAgdblxtqKdBp37jntSXPpiH7d1zsnPNzvO
G0rIavWiFLS6ykVun+4q20wq9X0Nbmz110JR5t8sw3Nm2jZzv+Z5E38oa6NazfMaDIBGB5beFykt
zhZynsIHnDONM+a2SsFx0CPTOMvjpwTd3+WHHNHJaRiMJcwAp7InB35VHqXrFih2GuwYpD6+6OoO
dWcomNYoLrqPeslh0Rs9hep/V9UWjk+gDrZsY0u5pTOw6PqHWZNhtcW+1ZXYAhniKx3bzFa+wh6w
EwVqp4Y/5fUcOPuyKVIebkSfFbp2E3dHSbIXXNPZOvqW6EqP1Zd2uVfw4LmNe1MzycNp49U4e10C
8GdIis7JGRDoMgExZysDg9v9Z7mT6Q+xy5Pb01wK+TmfCSyW+b9F/MJuNGArEekoyEu/g67fduA0
8UR+deX3TR6w+LTwlbbC1GkIefJejGPstabNBCJke9HNI+Pr2jG49iV8eKmuQAyN6sfQGhIZkneb
hidQw1g5lJHGHGp1l99m7/9rnXHIR8AS6P0KWlz7DN1SNPewVf3C+WXWV5ipdA0BVzFyOnndOG/m
tRPFYDLVrD2EzCXSFqEuEqGLchcjDjxltm6ST95Vs7amUqUMtcIPSzzKnopdrb4F9/T0k7dDgEWc
yPObZPOf/5VPBVKsmwGuwOcSg7NmMw2P/LIf5giW27ejDWY2FhIosI3wCx6JtWjecnPNuQOaGAGh
UZqXDKB/VDaO2b2srf5tU1RCxmsqGD3OJrpG8z3P7hLYrELjw0gphM6x5RR+f2OnOgzWRUJKvwSY
2Ocrb6Dzb0tnl2mfGKflLEzbR0qcRyXu+enTvJltzv9DjBhX+cWhIKDhWx8QwXQ+phm/O8YMYeEH
m+jJl4y0nGnAkyvCxy4fcxuyPBSWzRkYi+qEn//jqsVLOEKIdpQv/bQzLd/HjBBBKO/g96MY2JUr
/lmVvkrVdJsTfGo6eB43RTQOVAOW+Ms+heIPDgZqaXi5jLdWgzsrW9uJXBJ0S1jZ8VfjKSw6MHpZ
CwoiiL7IizvwfDdBYDa75aZPOZwd7Tn5a8iLL53HoCWJHphmH10+9e062bYmRue1PHklosDygV9i
pjTYW0vcQ6kcWNbyWA9Zvf5YljyUSbRkT/f0F4my6ZwtaQ5clQ6Z44CbXZAwf1XXkwGrsJgvxaGn
eCsuk62/Ypgvkdh9EyCpZ9dI+9nAInMtF0x9XG/3we4q/SxrsjCpZ8ousvRxuXr2M9QQ5eRouOn/
IS7UcYDENMuqSdGnB+gixmk/KDpnC+V64faW9Tsn+krg6MF2AkLcHY+OUIpBIwaVXog/9PwrGrlY
fQs09z78wo+AJMlJ+fdjL0PIr962bzpKGn3HTX5U4Od+CECfMSQocRHGO+dMoo3QZ9mrVP1ThpWj
8wiPYX6pZd360+NZWdyFYi+g0KOd6Z1/BoCpeztbq9SnIRJ8Dp2Wxk9xqO5D/XSvsrl/D55DRFDl
qi5kzi+5GXwHmeQHAl8ZeKhHwGdzacSgpj8tdAjtwZb1a7tN267F8we9RkgcWuH4EBiO0Z8lW+Kc
kOsqxtWX6uVmKJ6Tu8kixZNizxUYp3r9e/29pCRb4AznoGkb505lg2TNrhNPXxpHWz9PZnVLLY+H
ZusttvSUR3bK7jWcw2lE8qK1Sjqpk5QUlFNXsy+gXrB9z0MN6SwI++WkZIru7GM0nQ7IqvG+wGfz
YoX1ZtP8Mo0YvXevFoEwKwz8O7XaGJSHw2TQHr9mtyMLKiDEyhAS4Dyqjl7IQPw6hZwxLTVzmAO2
q4wma4Cn73dtcaznCAZRA8puCXqHHVT18L3s4JcBdsxYw1Qa35yFNGgbaJR0QMDvGO1qwE+X+siX
+vN6ede0ai9tZbhjo/XyCGDiZpHICTbI7aM1QWPHUeT9daQOM4i6Ph0bbYog6R2KxIyEpqbFoGXD
LJFXGgWp35thQhVyWGjCEMLdc10lMXany+Pf+JL0EEVXfhC5Dpcq0aa3d/dKSz0lblWVEOfKX1si
K54Sy2BUR1uSIlBwEiXReoev+rtofiNHIzpy5tIgK4i500VTCyl3KRFonBM8rZ8ocIHQNv1OOvx9
bRhzXor37YYptqJX7iyKvfPjzYPYJKvjWWmfLNpn61eJIgns/dtL2+u1I8631HN5rAvSO7tPmk/L
w0HJlQtQSxq3Zj3diVKEVbaNDLXORvqOixVabTEQY2tNIdE+snN8x8fiM3WWGC+azLgjL7VaCSev
WJYJjOaD+o4vpkHF4gdzW4d6Nv46AIERcvhzdAUe4gMDLzXSBRZ5y/O2Yd4amkcinbqqVrchpRM3
o3H9LyQBnB3D1V1uaGxzABfzhBAf+SDa2Q7Hq8zTiO44mW+VugrjppxIqQL437mUMMAWiJvXeVRZ
fyd+fa9dwCMcJmZytMZw7iK58cqorX80tUbmndFX/Un08cJPluh9FfDJAXbLi+4R9Snjm9FqGeIw
+poOufBHOii8GjIAiMQatdQ6Ndws+51xMLsFex9ItahKWWZ6IJU4dGmX7c5usUuWmpd70RjcQvyT
Jtg1q1lLtx+E5xgFV9eeJLfZh6lNmaUKjNWJU5x+hh4TH1uQaRdUmMPr6DgTIRB4gYg2xVVmn8rC
pjCk2FKpOXoLvUZ69if8ebiUGRpOLivh/LDyJgQBkLEgCiK7GEiPuxXK5dev/k+stc+DUK+W39ut
DAHUk65ffbhZH1OdTLemjC4c86ASTxcgBoeozzLDXd4z53tZ92i/2vsEL8J2DsIaEpGz9C1Ss0Py
yLdyIdKaaPZ6iiY7GrsQsiMHFrjvsIw8OyWDeATIXNpEenKaRxG+x9ZFyRBgxB+eua8KZiC5PqBO
N4/d5U9BCbNORKeLRVXrElpj2Xd7/XWWhG9e8fqUik8BgA/M9CUno2qR6ChOUppEyJ1E/xSipC6f
h3bNbNyL4HOQRB+f5tRgpL6MB6kccv76srCVawczK7SoB843hG4jEQ0dPiK4M3jXuF/Zh9EsWqYT
majeEPtQWIKLIrRPg73dWlYY+siIx88gehzIcITFFWPzNT/RPQamfuxkf9JdhI0LS3laqcYmfe8f
NezEJUguyr2rBVBQpNPwgN2QT1tQwCozHcyHsDbkluS/yQJHvpe+xeUZ1spEaR9MKqCN21xxgV41
INIEHfmVcNjc5YxKtgB0HxKdW8Rw2INOkTC1JK5sWTyk/5vTrBoFySxSxGMkBzdv7ozi7VHdYZK5
eCZMFUFGhikrmecide6dihWHynCMSsKs3Qqq0CUqmfbJq5zCJNUHg5SYqlpi/2DRdkjdVCxBxp5c
e2SsBzd9Z83ESuhkez26b4ndFqe4uB/K7nukzMr14eIg/1wgb3DYKd32DTCTTN32pm3h9WWMkd21
R56CzojJPQ8vvDTq8ARUrjTqXyYOp/aSbZKmcH/05TOpbVb71X1csUNU+UpjwB/SUB/Urp+YVbSs
to9G4NLTtzkDGPgQpYhFsvlf9kc5N+N64X1+bRmzBx4DSaOrHAuQR+I7EY1W9EA/O+Eoy5zEX2cn
wc0VIhLhArk/yxEsjUkk5ggrIEMgRkEhs8O0Oa1HYk3+uI3i3r9ifsl79mRMbos59iz5dfeUYxoa
nUIvadbkjAxD33WcuZQFJ6qh9LuNizwJCq+j30uSKLxNgy6hziH3NRDo4cn0KzN4ecO8m1AMKIoy
WjfxseLWjD8w7Rk3xpT3Tz1oNUOosm7q8AUcT3skwkWg2dSk4R8N5Ah79ha0eF2WujlKZ3tUylYP
24hkEuJ7lfswY065XnRlDW1cd0QDiSHI3eB9oyutoM6PJLKiwLGrjKKwwQrVCIpMNpZEFZrZxdRf
wv2u1gPMAyRwcIUTqWT/Qqg6twVcKWPfyGngHsk5PefzgU87sz2IjrDtMOC7xASM7l+yxHeiwiBS
Zpt5OxId3JWFgRRVB03QirNr8F12YfgzwxaBNMOHp1dnGFht/8KqCl2btZGfb+XPwgrVkyFMSIo7
58eCLOPX9vZoNG6EOcqUZzLnhNz2or1vY+trjadce/JrtI8n9P1AUhBzMWByRDpRw/4741D9zv8b
PUVKcPjXTAZZif85JNQU5tsH8bWejNCUc826P1WArVx0cxkgIuFDwEOQbGHwp5u6VRIYOpkjnE7O
hVmoiWKGWgQ4LzPSWNiVqTyPQ1BkJE9JFpKuHiXZB9ZOCR0YZYnCBLqaXWrn1SLvs+uTiCk9kaXQ
vEymGcMWm6qCBHpm59i0SPMfriX9V/I6tZ/5NzgP81eKFQHuo02bPzpG8zdNLq4GO2g7VrjqeaZF
Dc13TpzHT/ddQJ4bDAu0b6haEyl6RMHykUsdFIJnZ1XrXndi3LoGq0FG3p6WcgNdQxcgrTshW5fz
y2QhVd2ePS36RqA+yHIlBRSjFkR3qK00W2rlU0YTlDFRQ/Wqdy9+kTwIaqSKNnFMg8XwOvI3l7A6
ipT9AQtzUk0XXtTJnIBWq4huExXYLl9Ul4dWjuvYktCAIuxHY7YKO1a+uPn2pGj3Vlp5Cg36n86T
qMOH4qCNUW54MeN8ahaDNJEEIk1YHEQqFtXhMzuRRoJj5aZytm9g5PmCnZRALRneGpBhOBc1MgFi
bVFF7itwvi9gunJXZPTGj8t0aBywH3OhEp+C6l9wHXTA2ib1Q/lqtrOirkUYl5n3ugfoAXAMjZk0
3bPKrbDy1GTeMdO17NpVrivIFpmHaFnDdWTdnPyVGDQ8GIHyNp2fLivhYlaTSDiZxlcqlXIr4mh9
CkVyf9Mml1YAl7TrZDLM0X9/OQa3rX95j3o2doEDD6d6EV/gDUWTC95SoRXnRmq5gP5g9nv+uIF9
xQkrQEo2lcqqvZ9AMozTpYRUuX5HqsVTT0Q0SAxFPXj5D74m42h5k7G4+Yn+S8pJfBC84jhexrrB
lCr9AryTfGY3KIL7QZIYaKPkmLgXYcFtJYwPQHi4rYrcCpZ/4C661lzpEsLMivMqOAXIXB/skwBa
UWoPK5Oiot1eN0rKBdCExM2ObY9NC8OO7K9R3m1bq8iq9+2JvBFkIMbaOXsImSFXWTf269ZMXRNO
oZxJqF5nXsHaHGaZW0OzbxhSmitwECe+t5gWvghKIflso/FAfEJxepXa+4nGgtWMsh4e+ri7Rx4o
2EN/LRYV6bRu6l/oCKDQgsl0EJlPYEUY2CNWIn1wXDqTx1cT8it3mQOGH/U171DgVI70aGgp9a1g
FX6EQV1O1IZ2ZCwc/pnflCJ0AyTEnW7XzSuLZLR9mlSaPW1vgIfttufs7kNSQRX6F8XgEuczZW0y
clnZnIose8BDbGPNV7fYWmZ71JpkbOOEYsGjLjx/juHPDdeHmF3b/6VgUIc8JT8Cn0wHT34u5glQ
aJFUt38Xf1tw5TVhMBXSacme17OZpdP1zbmm7MndYVneYPUghLWFJdzHtQpDFHGcpLAvOrtuYbHb
6ACNfCmJ3fqy5Q0c3t/GAQIb8qY9WECvh/QFJtLC0TV3S/LF6WRtkd1dkzFDc5Hx3G4Wzv0ZT+TM
tZu3kF90quZexs69howcOv0vZv6W2YqSLAwLcA4tWtfb0+ZceUr1uaV0BRH2JASME4inV6v7KiM8
mSYXMaNQiCAzoU7XH7FtEiai2NgLo4ia4rLkCFAldBnVqbQiSAKgzEiKlptgaWza6WRz3+3s37Z7
j1axZveBjOuDFAlbRKgfFNWLT5aiuh+pViFugPnmsLB+X+o3gSbcSuu7ECbf6zV70AUN/bsdVDiC
VKK4k4tTMSqrHppcpcX3KwmgAsdlNneoTzm+9eQJfeOFyvh6ycz3w26K7QejL2osL5V1QCAtMX3Q
9bhENzVTQMlbSCWMEZ1OzoTcaNcxB+skJZzyhKbKlJQg9ghFr67HTPXWNY3RefRtQK+eonfldIQG
LXlacDUI7lnsgIzVOAyABSAOFCmXRglzzMHuJxrMKkNTnLzgPyHv/roTNFpg3PeB+1fBpTnqe70T
gikMpESCzljxGlBahwlb+tLli4HzCKs1H/NmSIpfYu7XLB1Ek6EqdDDivq11aKDmWut7W17zWogD
yAIezhFs13U2lId8jLFN8gtdn1PoR7xFxY9/W1EocTCfY7hZhhmOOke2uzYXMKeYzPCnRfU31n/G
0IftcrSRUD4IR53ThnL3LDRWVCZbkb6MBhSEM3gS0fC+BizhgOp2wJ0iPgUKKuLxoiSwkd4gn6kh
k60Xver+m/NWEGkLgrwvpndOKfQAlqQ4tHMmbxFnkydg6ABfy3/uVMUZ7obqs22s1qxoWYgrt3tm
94ZcjN7yKiTWVk7jbz8oDwiNPln0Z2VmFUFlUQiGgLqCDdHLtKIvd3CdujF3w+n/5Otz2p1471tK
W7S4xqya4v1U7FSeopKXUqPoboxQ2ot0Zm4DWUGd85hEhphDT0DZPbqqHEM0X/a8tLroJxbIasVr
v73+/wNTD+hM6VWmO6AbOuaf/9ZqiPRZuarUFsWkTrTGiWoHkj9D1Xe6jgc6MJYFALADohFNw3J9
GwNYr4tLcGa8Ygyxm3uBKlnaI9N0XJQbnv85XG/ZyyVJPDrUcdIMuqdEcQuQX7QzIOWl4guR7Rw9
olRo+NMMbQ3zu2jwJBut+XUx2irJj5yZzk1FkGA479QVvVoDI1FLUJFGvCmmH+wMBbpXfvcuVNTG
06MMLivWU492gQlWTa0tCVjgrB8eIMI9pQifpjjKWnO2HdZTfUdSiyJSGouJgKyZRuDtfEbflc+0
w0gKMMtUgRDwg0Cf7dElcCMCVsWOQdPRMdvhalBDfSA6/U/GbsIS1RK9GB4ZG12s3xDnN6F1aU8r
6hOyHD8o9h17pKqQc43vCfyuf9z+eVw1P3OAbDChy4Ko1VXMWIpxEOvdTup74zZ+a3F/cvSnUKHP
ndppjpVT54+5FcPoygsE14Q+kwSI/gbqFiC9lA9sxW3sLEQaO41eX6NUqCNMSdX5vp4iqXeVjHKH
e0+8/XYwZW+4+1HqEvsNYy+54TYJNQsU6K+ETiTsmORGMocImBkaj5fh7L6/OYY0b1AFJSfWG28Z
gDYQnF3ZipC4iEFecqbeenwV7KjNsnxe2dNOqT0HEh+EPd7vyHYW1Shm2oeB/8nTT2CMxnXCCxfR
HmnVtsyZcyd4r+Ivzjd/VevAkO1Vca7bFuk5J4qZq5Ysb7OTJU9cjvTG8O+RJfD8+pAQGdCJ09rN
/Oqe9fu5+jGiarAowCmUkJbNRJ24L9Pd0Tf08EpylGD8LyhZN9W6/3RKdLyhvW7DgocCJTBGE6db
TORcep4CFBL6eORC30rvjpetgRW35zDMb5WrgPc0BsAiP1aOoi5bA3p0AgAZcdt3lVqx/YeKp2rb
7VNhlV7FC/yei4quqgvrPtp8opxo3e0yPI0pQ7dL+b6ASLCRoDA+O7YvK2noM6UmPFz9BPtNAXwB
Zld/tt3SgilqhxepLgH3VG9T7NgF1kJBNe3diu4CnJxX5dx9KIwNRcnkLKObuE+fWj9B/5fE/SUZ
5ZlAdXccuTLSDHGVxuH2EW9yhqLmg3zoxJIbM2NKUxIID5sSTzaCmskQT74QeD0rhg4OXp58Ptf0
64scNk8BxUP043QbYaB/koXml9FsvP3Sn4HfQLpn6WsWGP6qBQOdjcSDQCg6Uk2w1gL4q705b/UG
AG/Scee/0R9+aCf2XQWCpQkTeqT/2HHeAa2+P9wYxIBWa/18GVpy66qpqAab1yw1pkIsAjTB3jZ5
HNimxystVHHeEqsMnVQ6JMouKJlystFKqwp8SZYaqI/BAuHIBxcghA/bS03OBn1VvHi1Lnx4mPT4
K9ylMw8r43ceynjgwXideQIV1Vvp8gJ6MY+LIMIsT0/mzP3dDXDbYJuhI3So9ZQDCPKclS4qk2vM
1tu/XAuXRWeg0FWkmyq7lefITaKP6ItM5C4EuA+yjjeAsrNpC5zaPoi6/E68fREwuT02UZzhpRjL
XjKrfzqvF6S5HSA9RPvmqX2Q+p7YyLmHUNk56HWyQ2BfzRCAFR35L6daDUPa0YaWDQ4AzhoIOsZ7
KdJwWwrgoFzZF+00ebQ3Mk1PyzOFX66fvUTCliqklyXrL4GG0mT9AXxop5O/dLOGZ3nT9JNf0kEy
ALWC7eAXUe81zy1LWqNkemKrI2iEdk7DDIxwJjkgyyI8e+paFzorGF48d3CnfC9WRzCkw/fHkEmU
wrRWM0MO3VNiIXD2f1gYkIh43GCkV84YGn7bD0z8jD6ijVjP92MyC59VOqPytN9zGPwjkqAhLPCx
5gDr/K/1Y3gCtxFktSqg/B7C1S+e4iw9ids3ucWDkpaIfMTI8TFo/QO0mzSSvp3aM2oAnN70qMky
OGwkLo6rTswb9BXxTrPiRSoqzq849//pGXDHYoatVvbzrxZWBBQLit59boJ+GeGK3BAoNKUCtC4h
6jRaaBn+2bGpP/wi7h88bEEwV4ytuQSKsTPX9B5e4b4CZUILk7gExAcakG/9voXwOWLSDGDHL4fK
XFPTvxGbAVGusXY55x9Ae3+aqLQj5eyAddfn0FF3Gqx84LwB97+aZXhjTxCTmyC9wYB9/UWZUkin
DGNkx+mC1rKdxMbAwWW7CvciU0+qtPYLvNuZyrHt3+MTaZFeu/np/fYwwewuFcfEo389nHbhZbDF
ROtPjdCMZPg2BSYSJB4zkMwgFHTwed/73SyAlBacOfI7botKG7sBfIQfRa/Lye8+442Y7MFl2L0+
jQpksr2Q7PZE7qLjk61TjKtIOYoUwFRqH8cnZw22AQ1qX1/9qs2ZpZsH6irmYcEM623m5yKSBQdb
PxT0+Eq9uTCm2wbPKGKJkqaIpLgSwk35+tZUGa+8OpgBckVVO+uL88RaMRUJkzEU8lUdBjC+6saW
2aOvhvO30uApfeadoylU0asJG7lSXoO+WBR8p12zgSyGch6UiGM1xJRgegkWYD+xVIxY7O2eI/1q
QM9PVVJFxHGfmthCftV5hg3Ot4l2rYbEc9sm/sJYI2xyNxsXdFUjv9rf84fEkVQZaXSOX8L3MHvC
aZ/dltFrfWS0VGDs8tpSoU+34vB+ovs9F5/MZvMsMhYdSP+SoWv92MuyuDvQEA1HXXqc8WCoSvGJ
qlOioJLfnwe8qkoA/mql16Gp0Q3WGMxA+YOFxG/nXcIpnYyFDapiWuUn3WuedTzxOvkkq5GqmiJn
ZbWAAnA33UpJ4ifryu13vklrQVvLnUmxn1Z+uCWlODKMSkt4cQcIThF9upw7FncfqP1DxlZNkurA
/vL8MJWCI4E+T1zQR+x+1BiD99cKjAG1sy7h1B8uppuAluJAd5KZdQgqFy5YhqGKrWuRpaT2kljE
QYhVKPwisMAMBEP9RtBd0zMdZwt1moROd1KFtog9edB23kdYp8C6IR9xBfgnzAZD0ikkoLriNHCh
Xbg7ea+A5mr75vQKEkYOHDcgwcJ8P2H27v/w4evdlUV3xDlmvWbj49IX+xayiwDg4EqU/IFCG2zq
Pjr+UH0CR3ud084ngVKtXD8epfW+sEQM1WnEfesZGGIW4a0X0gp+zlpXXMUHZ3Kuky/CoNu9aD8+
xlZg1tYgXSEb1msqTVdGiIrmk6llgPiS5GaOtuf85QC88Kjm2menIA9vKfQXeHKHUZANI1Q7JCsY
sYfkK58ct/QKRsPk4kUiBI+U9qYpaUMtP1fJV6H7SXXF6lP3aSHQfogJ0sChWQv+BGM0JntoUpfY
xtUQykL++dbwZsxYDL9yh5JDzMTAWLDfU0YVv2R8SplkneWXNHi+2DDP/kTGqV9jn+DA/nmEDahV
Op4FaeXcqcJWTfAzVoOos4whSLDAT8+x0HN20UgCoW59l4dXg/+DvKThXytWgs+oAa+RvJ6YHR4l
64lyTi6d4RcAMAq/3dhQe2k/e5ZmmDwZpCMIIeRcaQS7++Ke2qV6K+74D8Z8cAX4Tkg9uqORK3bI
bGgkLRwbAltqwaHn+FwRqZFytGDN6x2xc/pVN2hK2dG5JuMVuUE1NLEd9vbirgBEmbsEGzVVt89E
ImDPSvs4/fEfY/RAaN5QdFZA2QG69H9apHPegbtFhqXNW5EhR4k2YmMmxN8XgHlDYelhEiWKfkGe
/ctkVAaZ+ey0cMXJWmJH3SRZzQ/gc3EG6DkDrsstL6/uEAAjY0Hlyl+DM7l/fW0hDeOOV4fshcq7
z6UsnktK4ebK7hCMgKICMHZAAhBIDCg1Rj6Urs6wFmTNrEQsXW6QFjdpXkWmheOnwyJYYzHQ7bqG
diX9ab53aFQHfifusHuxgcfHdaCp/yXUEZ4dF9uvAhXiJnh/Lbc2swii/vN4j+DbxfPnEzn7ibmI
lTztsay7x7Bsb9iiV0La70PYWJ6vNpUcxYcjwGnVt1MGaeBARQ9+E1a5FeEcHp4xG4ahZSdKMnAC
ExvgG7BHN3ZJm/4oGmwB1ZfY+Gw1/RS0xvvfHD0KZr8/bxIirzPFBT4lYXWbCPG6X3S/JGzWera8
f0Sog/tYeFkhB6l7wUywCoI4tXMm1RAfnV1+E4BJa2zOKJN+md+tqYXnUBI3Q8iYUsBElqvSTikV
fHSe0XFw8gpyf5RtwyaUuUpJbybXoSC83qEJlEHpoyUT6yVTHFgyjTUEVMleQHP3yjcdTyegbzH1
HsMdfAFRZJBq2AJ/dVpX2KUm7RIP1MCOdCa+JwXQgyC8lqt7zymgBd3y9YM6Yg8ueqAojewgwYdj
zYclnxcW8b1nHstgV6vMaoAyZ0bxO+VMivlwDqxhfrxCZjk1Y/v6t0u8NwPLsv5KEoup9ae8TM1d
c/MocyNTJt6RcVBsN+TeLSMmN3ZX6ix6A5Q88eFjBaqqe/DP6joFiVID/zOoewwLknrSIf4RZPdb
zvOggdVdgLLrpXXku3ADEpOZSFf7mWpaFCCT+gjfQ7q6ZdwbOy5M5UAVdPl09/oajtMxERmoKea4
OiXouusfoFTV3szdJrYi8waA1s20LMzIVRjZir1KwLN5FClpMIvKh7egmy3lJpDAy09KcdXyYoEl
dcyW9gK2TWKWxWdC+6adAnpYet8r+ZxOyHpHj/V2R+sgKUUtWfD4Of20Gj+LGWgoTqSshuQ3DpHw
+PVcw7cuaoVMsYQ/G3FqN8MSUU6vf4SPVxHHRVstQofFKWikVNWSnILhaVY/qRKkhai7tMwVdmRt
m4ELnDQUwBfjf6oczmv8Tyx3ZVPsKePsb1/IdmQlaHh8ZgeX5dNFGJMfmW5H169gRm17F6Zk+Peh
VecPhLvkKAkm6RIP3pmalJAi8TsmaspMnA8nH4ZmqN7hNbMs/RjYSLeiqLzhV36FiDYM12198Y2p
XwmUblM14u6UQZ2kTDtUYZyPyNFJtad5cOdN1SGPINw71Rn20Et0bxAP3jvEJoCSA6Sgzjsb3STd
becr4b3jKVPyji7MpArCRcvCgfg9tBWCPt8Ouwi4wiXid/hCu/qT+TiaUoVXXtYyJCiKJ5GJtnsm
PticR3RWSprBW/hC2TzkyKVmqSLB8Z3cAzevIBT7OZIzmk1J6sPruOIXLAN6yXRrsgWZdvshZOIk
7zLWFfMkPM9C0o9pcivrd8QaZIKVsrOHtywoz0vtxVcZbAIUWaDozM3lRqYPVFNusUgSzdFqLorG
blqLKxZaWO/EeEux7kVlxmdxJlgAvG1PjEUolvBaaqWkE6aEGCTB6ZFwd6i1YIkwtm8/rhZml9De
PCDxx+B+jKAc3QlejFUP6GdQHLIMXVNvqd4YrmKXeU9YuuuHRIS0OHQ7UmzoBbBq7IgEFX3lC2Y0
ixXZiII1PP+GNO6YLJgqVb34WsMOUtpd1zrY0qudMGL9H/HbKAmbqeCAVCyvuHwbvL9Ht63MX6+m
aZQGCMGqu1zZgfqZHRQIl3oqHqyuVfKTKjGfOk/fMCHsSLVmYpUwdxQz1zLD5sE3Rq+YsqCfl4bs
MYTlawJF6PmwA4enZl8TMXLpsLn64e+J9EIGP8EPArp6ww8bslgkw0qrdoj0cXKvCo4734Ogry1j
evK1rnyQkWCaOd3uJWObJU6Wx1yI9NFwcIRJhD/Sp8iGR+gT3DIwHAC4NVrPelo7SN5R07aFyvlj
JcUpjV+M0f6lcQrAeqNqFVVKZH0d9k7Q+smHVkjV/iYvlufyZvKraaCFQm8ukbgOWsV6x4hM4DxD
M1BBu72Lkv3QrzqPAunX1fGR/M683Vf/Y+R2BreikPjZ6DVU9WljWDek40Nr1135kSQqPQDKMYnD
NMPNlZYuQ+EnVZZc3xN0mjGH3K7seo98Q5x/LVu8/hbZhZjLY2+Nr9dzEhTTxpaHp3CayI56GMjs
vArfUxXqzStb14pSENkmR2+17efnqRnzy0kkEO+DyRb/lJhP+UGqPlZIKhHlriOXwTnzxv8IF3I9
v7Z1AaqG34jvjVIftuvcK3AHV9HcXV1be+Ixl+gmQLHwYhsPRMmgnuj0ZwTA4b4v70efR0lqljoS
HqEMecao/30teo+xepUVuj6shqhU2J+7enABjr6vB1Pto+WbHnM5rnLlRH70VOFumNfMJL0nkhtn
bOovHXAdCy0IFIe/uLX0bl0s82w03oVFfW9d5rcE2LATlKBBCcDtWQrIcDI81q3kNUFLRMfeqxQl
6hN7qzCd0Y3q9XcwudjAXxvYKOnEOI3yomXbkwTn59ddZB2hPQjbYXGmVSLFkJ4bVl9p76C1HQgp
PmcWHJ1AYjUEgpSAhsrB18/J3oigaZLD+yjMkoXKTKH1oAJbUIdFoFrIPwpsZECbMpgFeBIt/scW
q6+sfWEdDRjRYg58ZvptS2HL2rO9dIY6oC40/r9KabDMmgRyv7Jjl37Nm+tOZNFVzFA5RkIg5W3Z
NFR3dAIgT6kzsouvWjfeOqCbvIo8Hid8kMlObsaOEX/J/ceJZDNmxIB+B26DLWCik+Yay9lV6iBR
dRIXZh3qOyHmtGZ5iW9umAlC2iWvz1HY/aXZ08gZIt+0sJhzWvX9eVX7njxnBUnlkcy0eYrNa16i
9FxH9OSgX2ZgPPoAEE3PF5WcuIRWlKpzv5bzG01RoZ3MK6JDVn35ZVSV+NY8vV72g1BFesyPASvb
SAEMH3Hqgc8bz0Gcqe+oFPG0bGY+t+35T96+5RvppT4b02+ASTMTnzIXNltfSkZvtgWt1MeRLpuT
javZnD1PQwGpwfPVE59GGkeRzDVugcZzD6aRlYF7pMhSnLPQ/c1t5znQ+V8HRJ5zD/O+LFQI+y3q
rnSxnv2tBHlS6azt+01cfO2rQ1XuCWCqm4gnmGkN9//SpiprkcBuWpsKECq1KorieRrRmOtOCgQ0
+sadLNQ3pI8kJ8MvGN6BBhKKMFtp+xSDlcntdyb3CREBA40V1918idpzj/ZhYJUSLlJObyVcX1oK
jZ/1KTyLAOniPhHITpJdvvTE8FJ+FmCAxEhmy8u0k3D0cdb1jQMi+FGpxM/p2kimOrRrfq2ut7qx
2KFiUpzRMQDZgKSZWt0e9jwdSLp6XnV3APi196uBNNiBAdIdnsuwMvcHtjieUx27BWwPevyHl0b2
8SSFjsJoCPL8kxomae5ks5jEEsOe1QONrb1W+aKRHuj3UClsF30XEPDM1BushUblHPmm9wum7mQC
VjXYvl9I1hsvVXkiv8UiSEBpGc+o3hZPW97BnU3YVh8PCoWapXHQd4IHvpSlfJmvlxK+MNvxvkpK
H/nB+y3FgWtW7PruUUu7EQIF59jKzhf52UA5n8dLQA/yIrbb5TLKD9Fnf5b5NP3zfNyKzGwiOjUW
hUqOuMW7u7TzMaCCu038N3kBcrS4END6CIb0Bp7kmUS+9cbeJ9SL9ARWG9myqRMkGj67svVY6Ktc
WklDMVlmMvnczhvwDN50EIQg5I9tarRJIfKUZydYVBPZZqL+OphatCb5RykF9jxmx4+1U6myoriw
CueNiEUrRekZ2hcbBAR1JVSAxEERDlR+6/YyU92VtFSt5ANVygZ3cBs40Yrq5MAwUOfQS8V2kJsG
jHuw0WugL/S1U8o4UXDVJQpomPD0G/5f6QEx/9NYRSvsmVOt8anQN7u+ptnDT4C+T7Fb+QglBBXV
puuPM6wY6gznEaHY/DpAS1m8cskfWB/u2EhNNCKodMWAjfoOSI+CtEarrqf4OjpSIcurtvtmk0AV
4DP3Dsl/1CYNcVyDi0vN7TDWdsHnqqYiKIbayizppvXYZH9eeHB5zaWgtlEyhq9ekE5g+WnXt86Q
XXwN2dctwG4cozoy3M9ymPwDZoc34Kk7BRMkdB1PZ639+Yupx5jIAEZsi9FOF+XW2EcXk2AJdGZf
n1gReYcC8INLmFskEVjkwKJt/BNXR4+7DU/h5i6pONN5RRMEyuQFViYifPzNxgw9BT8m+MBToOSY
0Ezdj28o9FSz3blF0bBzLDwUcCiExq9i9hIoQncNPX1QX1cHRJt5hJa67ZrlnOkAaaZHpl0l+GzR
ONFglZWgTDPZhWfOOUH7vbnSptgWxWXOc67Poce64/g8GC79B4vee6GLm4eS5vZ41LIpLzeWyBV+
UBooRTkC+YDny6+9MjlCQFoQ4ZF0dybp3dCFy6pV2VlcdYv7UNv7WNq2vXhSLxl0Qs9GvUtcdToi
a6HZBwvoi503/eMwaq2eDTJ+V73h80ilAde/dlY9gQ9mVT5fMKl+tNe5mQYpyntcUTNwI8EUXUuz
LdnsFO4fysbzvfzd6raY0LOweRZk4FE/RQ1iCGgE2Y2c15zdxF5BWY9si8OhJtPKktUK16vGtS/p
+T/Y+DNoCXg1M91J0A1Y0Vr4Brq1cTApXKPVgGsD7/Mb1X48KB4HOMBYCiEAUa9FSgOacVYx6DeF
Y+ynenriDxLBh3AkdtCJ+9t5pNJiGLPrFgZGE72h0nvdhLft0RHOJqu4bBpRC3TZ0SbZ6VFK2BjY
mMGu1LzBhFSXjcSofYOphrrcf1+Vsp1IpMf76Y4pYMTV40kkH0ZvmBbklG2XnqrDi6pnnew5pto5
6ANrVgRVq1O/1YSMjtcIeX11JzndsHt0R7yk0Xn7NHNQKLEQIX/9RZW7cZqo+w5OTaf1FFtTZ30I
AZHigI8Zzm977HVA3SbXibQmAnMokXi0xkH3lZehGGm7v1joJ9hESIP8yxnqwdHq9qk4256PA/B6
5ZYa2mKIRzolWXPkRl8Zq5oywK7JBCM+XBrOBgK5exoYuDBkysZHgnUgJpL9Q943L3uFZfUuPyMY
4HVLuCY2y8zTYyovU1k7TcHpxF5iMR96INRBAEoCDREdl0G00tA05ByQ7ObmFp8LlzgDhbTtfi86
+ZH7JmE1kTo2n3+4un75THEDWeOQlQF3iP4VG6QHx5PmyOkf7GL0XZoZTh9lS9Yt7QNj/oE2vfIY
tYRqVlFI9fwuYPYruXsW39NdxPxeGSmOA7X/8Va8HT9oxQSDfhIHsO2e/boV9w4aeGK2QFNrVLgH
QbR5WCxQMZO2zTHiR3DjaV9z3yqXcUTn+m+TGnjKF3l2G/BbB1/THGXHnm6j9uSqrp+nS9R8U4dp
oTa+TNV5CXbYTV7RSaqsnny11gh6d4i1Hd+sZOJcgaYseN0dGGh5USS0Piv1TVPgGbw7vtpQ6acc
vCY3ccmPWnbXbFfH4Gkh+k/sRcWQDl/X6zG6hyHNgjZdGEQSprb8c/fZ0NumEAs6jAHTMwd4pXX0
fEF/IU5cri4IbeBxXYUl3P4q+P3YERAY0uqbi3bVb4ybbzcBxF1VdRrftbGAYBcK6fj04QUJ9ahf
CNip6q8qww9es5KcBAA4MI0X7xIT4pkl/jpmappTVp0wHqoxmoXdHYbnHTbhjdqhwkZfR5T2f1lO
QYBDpv3a+laVRqKMdZZEuWCq74gen6NLaeSckVQUejuAMoNXS+fwWhkioEbsa3YSh2VAWVY5MZAh
VJ343xqEOpFisD5eJ4RIYMLnGzZ/Vo0zQbk13Q0OOFWZ9UNiG2ubzRkXpuIbCLL4nQ9fd+V/V/Dy
Ca+M1pAeI3lUxV4OkeQmIcdFSMdBXsKK1sxrcMfc8BgBHgyiqYz9P4KKVI9l48Ml/oA9zcaviCgi
g7ad9F4T2rpQ0or5G5kaIjgPVCSfBxolzYhNQW/B4PRByhM8WURpj0tEj5DTjtQDrwgILlWeNQqm
RnQfPCfcgLZ1Uk348rYxXcHpPZCvTYlaeM/EKM9vLCvquYjeITL4MZkvO+1s0geSa9j55IVmiFyL
vA9qWYUu5PaSpbepQSsBWbkN2dF5Mr8eX8oF0JiljqJZg3HSHvOJpxSpfTVqaw8YcuCHNHXET6Ew
g9MwSdnpc+SWwWtV32hLmTr5pNdGHhixrfDfcRK0GqAWSbfNBKM8nfpmM1mJr9h0JamCUqkmxGin
GmLIA7oRROCqEFD+zLF4lrHU13ocoZ2uZxhhZ8pwmahXT6VDdwQTCJt579/7JwRjXdNMenjqKLKn
Qeht9NvWZZ/r/d7FcOtqFbMVPAJTb0TbPODjgVSNCPy6w+DLWvN/fn3EWTQZozAAw09Am9V0fvxr
Q/f5kB4HBS1UF9vgLsYyTeU5vgr0PqNHOVtjzN2JfbHjAlet7MrTCotPc04sE4e3MSUfokZpir2f
wOaN9oP3F4ZnWVR864lbavkiatlD5mrlea3mOnyq3kxAVDyKQnpVpW1I2l2Itl1IwI26bGGGYanC
PG/hPMWUZ19mQXCGyb105C537Wa6NwqftOX0YerhWsjZTW7v632tHY6NG4Aj139Dse+npXakhYB1
uztd+b1dPLPblCi3nC+dJOviCpVaRbsUlF3dfxkZvsQ+cRtZTN9pBguA/2O4YMq0bqI/7aaQ9UX/
G4xnU8Kiw4GIJgQtoiZ6ltNnAD+jo5WTJoFN96unOsYgSgNA48kRPEwo7ggDZUvvSq9+e5qcdQN0
B/E/tLTdLvPmamnqtZxS0k6VyTjq48cXJf1341lvHBMf7/BrcTEXsIa08SeT6udh/HazC7Z16aW4
9wkA9UX1xKUdYcVAwr71H6TX/EcsAd7+LAN/s5lQZqaCpu5W54Vx6nAz3gL/wqFfQ87VVWAvciIX
y7hWMFhtz9Q0bgjyFPjFKJQ4NsPqYZkBvAKfaPRJkSY8XxlgUnzT65Kze+VlrWThxd3ZZwPjRDR9
agTTJSMkSpRgaNwu0oY5t/xypik6bEJ5fHY8a+CK89RsKRDPTxx8aPo4kbZTFq+R26k80u7jG2Rz
zYpuGje5apHG3t9KIDpnvx+M9MWe4uL/mgDkQlUhFY6MqIC5SmkGh4LMGFEEviWb/zFxrDAAjWFa
iMw9FU3iAxmyIqidz+LLdelyOhuqVwhAWEQu1alzBzKLw3engneNmqzdcdT0jzL0fDMDSBxXBGZr
FEdTSdh91OMR0DvlyQ0yL0R8Au5RaSLdkJG5pT/CBErUSA7dK+0HuVsPrI6Mll3I1PXCZ3O1RnkG
OKdOpZI7N04MIZ+Z4Qu9lKrW9v3TDu4iAg8jgOffgJuenyBugqzKLNYQhgKIyRDPePzR/gJCctjS
KNbuBjddWCz9cTNTyTOqoFWDE8Km9EGi2i2Gfg/kZV/I1utjcNpWQCvMTTfrA3RYz4jAEM8aQIrH
n2p9Do8hMGfdVF3nSAm9D46qkGShpIVHKQ0Y3Hhy2m2khfZ9kRYcwL6dAkeCVO950IvLzTJzoNk6
igeeh5IhdyDDKxwXPlIR+P+Mpf+B/C6F/dbup4QdVUhl8zfMsBrHcbJMbCmzTDcRwtMWluTVHEMp
4ED7603WDLMUCYa8ovoMaDqKOTRVqZhBTzjajHkcmokdDNHIzEyI9n1M8Vn/kKgPHTbuB5to2T4w
ZmFY2R3Kpc7qW4EddiH0gtBhatzy5xhy62wHnSDRumekUIlnPb/vzPMg/Bk9zPNyMqaNZGB5VMFE
5afQvxjBloT9yUAYoifvq9pBRBrEN+s2vgygvDDuXZmZr+M/dpvz1GQYUFHrLNbQKtEAD8PKvzJ1
YVzOxqE7czxICIFvGePVdO4jLSUMBG9ikFHchMNPdLThmx+N9kpU6NR9Fii52lq+3jv8trEsAzIS
AzqWMHnecJxasSFQz+SB5OCtieO9DjTOw7nnv0sIr3WdhhMp7nrVIRJDE1trzzjWzHVEsE1ZBonI
/LDPkn5VPlgHPdTalURk7kkfWFLTptrt2//1cHTXYxuh9R3gVxUXjHGt3r6NSlpZ7pjmU+bb9oxB
EGMqFAWLzwtaHixek7u+3zg2SNb6KCZuTRoCv71MTC6ytECRHA7NtCM/oLCB862hfA8tWmqKHNEV
b/fNA6qv6azr6HpczJcikGPO/k8fgg0kAfSWgbHlcoJdwiSOVcy+cpOftsYhP1bmuLoY+x6d9hHg
NHjo6PogOLDcGcgH5HezinlhrmIQFcOeDYy6PlH9eRLQzxjEYoB7URDKK3K6i8he+W066M2ZFKKv
fgl+DSyF4ia6t178rMpjKEYYuNMn5LpjoVlKZq4Scgrxc06anCAODv0dTJdAB5KU7f9As8g5x4BL
tzalvnJCuw/DjLNBZXjQ91R/z4bky0ncVWtOEBmUujulxRNTPoGPsh88tPNvtcMzLtJ70vfSBPTR
UmHDjk6OiQET608wNhF/F4HLqP4XoBSGb6ASYJqtzph44fGb0TgOlMlkWJJ/xtkARkdNugblSmx9
Wnw9kFFlq3kM1NLRYG6W7EduslYYvcS6e2+D95i00uobUrWfH27p1qQnUnkB00NyLC96S7spQxpI
2kuqh/rm3ShaHyckh8/mqAZinFKyjo/6OB46pS7Mw6a2SNLLaXzGzRl0R6AaTnRiyX/kiMV3PgHC
XUFZwf2FksCF3NuoFgATQrgJNtoXsxJlQaAWt1AINFAy0+py0AOzm+FqoQ+hAUZ0vWoXCHWTn1zd
VFG397hg+4LgC2+Yo11gGWt0tlajqwmp6/kT6qrpaUPSKjj1WIVddYcq297Utjl0b1TAr9EyqSX5
nTBEVFuGlzRGyesngDIJqHlT8Fy3HRiPcowGdOWqhyQHzfI/q8eIMdaHmGS6CI1dswXLqRfSIw7s
Ok9MbDl2JrWXKq+IQzZ3jxZsrsf6bnG2hYwtAAiSpTcuOpDWlwWUOT/kWEz1MzM9ne9HlKAASmUA
/gMcWxIfi0pmRSHWaNVHLTKvadrT1DPMgNdjETI+9X886MKYn5tGhgM4/Knqs0PamaOGp9180Z7d
0Ukm5nLC+SxXY7lcm1Pv6Z0Z3U+8mQWBroaKlKssYDx91Eb9wS8eiJTC74pmTsvHvCFCkCelv3Vk
B6Vf0ZNdcWm6u7AELkMTay5Dr2mFcjWW7ue5HlY+WNCXwaYfT926bQD5FNHjB5ookr1cP89V+GTl
8Uz+0TW9nb5wVwSMkuama1Mr+KmLRdCd1QPRZZt9o78/4J2Fysax0ZwCZz0ZO+JbZGSR2FiYoO69
vDjW7kto7PLNGvCEvp+PGZ82QZIcqLCZkVXay8AaXLx1mNyG7KbcwuLqedjPqCjHhhktFJnnHT22
GqwgL4tots/qCB1pg0LAfPPYN3a+67/ccSvYwDA7OPcnAq96kPBPnnz4oMjYCRWHDoloYYXC62hH
XGzucz0eYgcbpJ64FnfBrv2CnvamLzYXiJuW0RAYRL4P2YEisgtwHVl2pFlvFWVzdYq8P8Ux0Xmo
/iHKoCOUE43zt43SfSs1tpwfuy1sGMe2vf5ShrMkccrOEi++z27LX3krinYZG8sw1z5evFgTCQr1
/4OoOlmsNBlHy8ULVcVGFSVnOTz0hBlIFaMz1oUOJpNeYCylQSl50n7YTKiGn1z65aWkvY6oRgQd
ayiM5A8vdBC3T0ahk4gVr8mGaSadRdsUnQhBVLVEsQMbLuQ1yevF59G7QEiefeoYf3linVe9rWJi
yMCt3+RN9j3/KtdQt7k+u2S5v/gr2400h660153SScgjOGolOegTdGtoomdvTTUqYMJLAURu0Qg6
CZC+at4Lcc696MkI7ZqnCB3xvNTnJ6pPaoHjc+Csyoq3CYoFBgHSNhI4mb7Z++mbIn9+eYlZboMe
W8vJBs4eUqMWCTRCpzIwtFHXkRUVZerdfIGsEFivez5vYvBlcyWw1Wyed412cW7aRoeWIIj5sq2v
o704ccRzBhcmdB6oujRGakRdzsVJ6voC5P3/oDAtcgs1gChINRXLHUbi6DvJ5IjqMCQAQUHYQwqJ
ufC5HvHBu6gytAQmKfWeF49e0GKbvKuQtvFwQ1fWwfvzNVDLYfekQZes3M/cEw73bYc15MnC5so9
uTLBnz1PLaDACf8UNqiTujgncFvfmmYeXREspZ9wuf3SGZfmpl3mgZm+SrZrRZv9sLZBaLyLYK0u
tL5ZXWG3MBuryMkLWetCP2IXR/o8lH3YWnZ/UqPWXnfuOnPufTMVuD9xHsbr2zkeEtnNKuyqGev4
C7VzCLdAV1QVK0ag+Thl2ijnkoVtu4KU/DmxN1bEqqPFd04qD3lfW2E2SF/kgHl/q3ihB7RxUrfy
Dkllj3UOvkCqHSIATeJxuUV1xZRUMs1BRDH9qwWStNs6ILl+dgGQsV8H22iV7QCxaKh7wbXCKi5x
DJc2tzCBNPFEpjjlNkhtmBYqwMFWciaaiCOjvQZBXT2+KzT/h+ljs2+Cby3B3EPJTRXrlw/5YibI
16POtYNJKJSzlupFPakAs0aj+3QnYiq63wVX/THpV+yq69TvCfkc+WZGCyGHsvpQOBN12dEvlecx
hgJtIf1Ks0kvFCOPD1EMHKhImNekUS8Lw4LXOzQQv4YBjdYo+i2+Kg0uMaybXkDA84yBoyBGrOO4
qXxs72S1bf7gN8pslp//E9QXarBgIRos7fdmHIq7I4AkCHpCSS0OvDoIo0jFG9ZX9KfL/G2YaAQV
5Dr/V5rSdzPY+C8B0BuDoYMq3q8P+Dc+paEDwX5uA3JvCm7Dv28zVJHkpfbGXtMFTvDQWZACmkIG
DyTbT1oaUAgE0TKoiW5qqWcNLYFsrLMZiEUxmKNNh37SteDd2Qmd5780sxDLylHunF8Wm7aqTf5e
PzrR7nvt9jVE72NvZL5THQpWWAvEz+yjOU756GUWIhdrzw5HRg2WVofdrTJiI3xqtGS8SIAD7aI1
ENbxCc7rn1sw4IRtieQIhoP/E5xQkFKpAivKmpZeAb7PjxBd4RJ3s8mrpgod8dS8ylWiY7jFQ/UB
eRDYraILLPmG6fzM1mB9rDQioIlAB69fMA0+B7gyxR5wEsxMbQ+hm4wM+bMZvTKY+P3IoqpMB0jx
xZg1B5xeVt8fi5xR2VyXd7bOpVJXwFdbYRBXKcsHHqLPZaOKr+CgyCYcvefwX9ENge2NAJ0kldvb
Bgjvxat0qo2G/FA+ZwcqNiW+YB+Id0meecaX1ANV2h4yPoQg2HVWGoFkkbD2zaF4ArPH6l1F2oou
vWCIzNj30hjxTmywwMBfZwYDHBNX5fxWej8Cl8BuqW62LMrlMMVabLNXr29LE14QaIz7+qaRM889
8VQE9zzELDPqaCcpDKdK/apcxSMTX6kOA29cigE7hQ51X2ysQJ2PAFueg6YS84OFx7Oep0pmG+88
9sgM4gB0S47NE4tSvqaWzVWW0thNmiWToV8wcwhiEM9q+eSdpJyvXkEWAas0cOgJWzlWR6yOQEND
7oRcsGw7GBs6wQGaieWW2w6ylAekaocuXOcxwfQBMNToOVi/kNMsPz/PFgkEhfk4XphY0CfWWg/x
exJa8ZU8lmwPMVTS+F+qGSVnqcb6k7SvdEGu6e9P6GeYpTN/6hQrMBUxnktmK22vNk4B8JjmKNTs
bIcC0zIo/5etI7KxTlbG2s9Y/pRgTuqGiDcXKvfnrJpWsBb7p4PrSfCqaQ62Dzd1OOaxjoRCNtZ0
Zku1FthZQbQg2W8m9y0nwhkaWOMmQ5L5tabpik/SgKO9GsCpi4ObzfF4Z2P2mx2mlelArYJnV7Kx
W1tPTPMXZFuZV21eEd92YrdBPILVamPAOkTLx9dfh+PxjoXU6tHb33yORPyFSaS1Gqf82JeCS8qF
YEbivKaJLiEzWGrmwXBkF1ecoNQpG542L7cjl72yDS53nHBujS1qFGK2bTZoM3vm/5TnmM7F3sXE
WpM45a9mjdRhnzr1XwQcpel50rSpxPd8cf+/LGOi1867gO7RqZ5X7G8HyPiwRbXj+QjftJrLBppW
VhzpLsHzkAofn42+pzJ4nu9cNdgukOGq18krTLkVaEMK0+eNwyVOVFpGMhkYxckLIZ+ZxDyxPXlg
t9TUXrQTdlsqouaESWRrXVkqouIwgZW9kEbpPiJH+eh4yG+zhDygdjnPaRsiBkdKzhk3MKjVTA3H
HuLlbJJ8MGhVdF+QpkVDrxttrSbiLUzASz14dFPitLOGpD8AV4f0udZG2BH2P6NuPVjwaR05hJTq
r7oF609cDqTkkjSdES+ioSKGUAgeMx2HfemIM+cZaHcJeXi2ZgLxKCnofzgOyCTTHZ10U2LWCElr
Ur7rN04NrvRpa4Cb9cGSkuChTHLDltMaWymMoAQxtYIa9Yc8r9L6M7JbD+x4yYb/z0YViKhtreqo
chLWOB7f8irMzERxd5CFkbUIkoGw7g88I04ysGUEmqZJeApcZWkhKR5nRmRm6X33NOVNj9E168kZ
l+hHdCoilx7LrGEaM2IxyUqkR3YYhEDylE965VyWgKqYxBRpqj2qRzWtjUHm4XKFX27rE2uNGs7B
3/dFHjLALEMNGDQX4WXSX0JiCTwAG5VFxjL4JSwagHXYvhJGDUhjDnN03/8++ckRQZ262R7v1mKa
mpSNfXD7mPZp921Pp9BpnabQTz96sm47rI/VCsvo0/iC2a1RpdwlD/pwPR4zXvR5++ageQOBPQtt
t6kvv+BAgAVNnc4+gHquP/v9/poybxS0MYykaGrsCUSM8tI45PeqhbnvtNz1CMp+8W+bj7bz6peH
8nbeJLYZfud65+xH/Mo0va+OlI1ZGJMaP0yVndirz42LuUB0fKd7c5Tr71mZQ+upsARZo6a5yXXf
ML3eoW5yP6QkgqVKVVq1F1Q8mhdIngBXpqltytk4eKKGqeH9E4O+3CuLbWoK8BQ1otKctvdhL77j
ZGm3AUpca5blzHu53JOFWyXSer+2JCSgiY6I1nEzBf2ZZfyn0I+5PkwGPIrP15Dg8ohcaLPYdO4g
BBW3HXKwrbeL8s1o8YGjCcuJIW9ZDXsNF4w3dAWju75wFh9iRZ/Cdw8GzFLvOeJbrTaRFV5w2Q3B
ql7UFa1GVXWE0hAInqKhOSVapGibzW/ZLQ9fac9w2Vj99/J9AvvSaXZcQpb+suF/+WR13svfRUvd
VrIoiQNUoYN4iMjXV3YUeq3OUkdNwBFfwLn3hMfp7Tys7cHNvH+JP4Z2rwJXASotOfLSEWVTGtri
aOC/5HVVAeGJh3VaeH1+3Y1R3qdqoVux4J26flyO+rKdP1BSr9B9h5Y6p/uMCEvj1gWu6cvlORSo
Tr2ismBvKu2EBtEYszaOa5KwQGcsFkGeX+p2uzHrGZg1Q9iJDxA9/WMFrad2ypsbaF9JpaEvAhlK
C2ekBRyQI9Aa0vhU9uk3BKZ4hWEIgnjLd7eXIDe3r0bNa7BjwWVWu6/Bm9LryUjl8+iHefGGt/ZL
oOKz8ZSUZsPOWgsBEICuKeZdRRwK252UVR2niaI3Y31vSU8lpjkZdS1gWtb347iq+DPiQqQyuo8W
h+bqFfkO3lEOeH7b/un6/tAbZ0zPZbyTYZcIJF2zsPTESQPdoGVkfLqmTI6X5aeqziud/guCHA8K
hXDqWS3b14Ux53L8FDv0gtf4t8wmQE+2aS85bCt3g9hnCyXCEiV8OT0CFc3CRonp422AJoxocp7j
AMImfPFfGKFLsv7BVQ6Euqz4pqhU+tzJvEHIOkMq6SrdStbAyNOORqA0lSgeqJTetb9SzLkxP7Xm
8c8UoFY2bz3t2QAfeksVlg7DlR7bcnDm5i4FJRKwPyOEQvI/X7tpOqTT9vnDVY2Ow+QzZFYbGk5u
UmHEMU3siSbmhJyTZ+5GvwWXf307SrnfRWuSlOxf62TRJN1gypRIERFA+nwMDU8GuA+FUX67/IH8
eJkOpwC9hSD7g53L1LYLTX9vZ9keMLmQzY6sXPEY+xVkdKygD0PYDcIFC7N54iHYbEBgD6bw/G8n
qNaQ7sRAN+ht0j6jolo4S9FZTKICNNFINM4Y8Ks5whtMhaJ4VcZll/coC/9lR9AirEDWZOBZarvi
sXEXU6CATMGY5mrN8Zot8kbAfYcum0EhJF1xltRWrgL6BiuJ4TOP+W9DsjsjvuGD7w0BzkIkIO9L
7xagATrq1Riq2mVOmhCsEp9acTjeMCqZK31SgSl3DykYtLzqVc7CxJ51wb/0T7cu84qLR6XdCtnY
gOs93k0R9pWWZnY5w0ClbYJB3wjD1iSW9eNVvM5vfFSFzqgWSR3RiUKv5lzRAaYW2C9jL2CpxCQX
c0jAjrVi7r2Yh7rLbjy/dbTmtA8Qb4OPWBGWOsPUsT5qXTQ1HoAV20AxPsbffDOuNucqZXn/douc
0CsUFAzqCLw+1kIf97x3MzDEWDNX0vL6YLftqwdprjOwfao4/Ldd/BclZvp9p/r4Df9XcdyuZw9f
C96yoKxl+MKP/3aSPybCGtDVsIHjZBNgDIEZT2R9/UAXDvjh2+i+xP7tUyywNNPrGZRfvJ+eobRg
qbHpXmfz6pPM/C4KllhdU+wqcu21xpp17QON8ZejiQvN2O6E9vXxO3AvMOMrvMPEjbTpawbo+a9S
0mu8SYbURHpJxm2vcyu7KSs4Nuxc73Vk7LDs5EGrGltn8x3O/uwCLWV4Zb8/jz9d+yDVdOjMjR7W
B3ZQtCFeYXlzrarHinYJycMz1R2DnEQIQt+5Jaenb90fV5n45PYlHeA03v94TUYNLml1Yd67Ynxw
7VzVs3eJABd0MvZolxtuK8vjUzrdoGTJ0opBdJkXmIbFxt3aJcUBtfNUZB+axO+Z4EvEQFnGc1Sf
wTHJH7GSKz6NQa6j4vbGl2Fi1wG4zWtgH0hWNzXb/xwQ8VTfWXQenWYlUyTxWejKpjvzw3gbbjd8
UONmhGbEm3x1++/Tfh+b8jftFx4ib5hQx4JqqKtJEPcjA8j9imyExm+bpmMRQukIwSpXp/3zHfa8
1khs2zDZrPIHp98w4v3yJZKJZ6k5nsrqTwGazAZjzeaIQ2N3VfSktTVz2aCiWORCTJ0cLou8RJr5
mO7VBwAKEmZQ/ljcMTPW0PiW4/ymS1XNsPXz0oM1FOB127UHPDpcJAO731A0COPvW9xA9FRVu4SK
y+6qxMTpewRNqzCZODR+n3wijTBDbXKaFhqFvED77Zs2+feMYRj71cHIdwOp9dlwl3Z/leLZI+H9
ppz2UnjiYsyIb9cdfbE9byUd3DZEPWojg5YOlXOyAK3JxsH0CFoWHBIc/UMWuWdn/OrLEOyuOGxz
rpCg88M//PgcI/AV+kFn1KOwoMcGblfQLZgfmb8q9XTtB0c8gAIVJz2WLSfGk3+Cid/tCU0egZoC
Z7n2dePcX1c6dtqvOwSL3EXLndhtllCR+xqjUJJYE/vU0Qm++VtUYwsKlY7/gscCMpKbevCyBu/G
rwwiStTka8OhM7Fl6jVyAmnWkmGviaKU/fzu+20JosicjezwM9ghEbAuAv0adpLzIaWLjEi/tx8s
y+pJBjugzT/260K0Wvt842cOtj7WGKhQe8wo0nlPSxFNZViCNvOxvRZyrWu7JpVkaPpnkLiyQiYt
Rg9zOB333kZ+77rxG+yLn8GO/PmBBn3TA8k5sBiQyY+g8EXJdqUCTBhIHw4x3m3G/fzWFc1W+UaJ
JRjVRTlfrpjcji6838ls8boTTiS1x5wVvoq5HsiWpgqEqPxRV89GDuAbKRkzxkVr4ixOXYgdAYF8
V2TG3yJowejcIuvGfbMgkklVAhVYfZaC1aX069Dgn68pcqFvGdlbIyLxSVoL79fM6ZhkIPCfVTqL
ogbdgfu99SdEJ6NT0Du2EtJn0ojowQvVRKVFXUZ2KqLAdDBkvsGkiAmC+T5x3KQ9sD41r/1cOfnm
vbFnFpRMTpRJ02Y1xdk5qvG/4M98jlH/4F0ehtYPVhHy44GYSrZI2D8oCiwv533EmQfHmEf6uU6i
61NEFZ1tCP2Etuned+AN7kFsOuLAKjvv5NZzEI/xjyaKO1blCTlWZPgMaMLGGdVZGzwvg2GLVKh7
Os64/OtOK6Mx4UYFJubRjbAZAzGKim1FT2xGGoW6HbzTc7DoWs3aR+FuQ/NxEZNsUCQmAupcvOau
keH1TcEzbE4mz7l9hDPqAqAXfnnL+R1R0KdTkLloAORQAtgWOKkY7/t4veJ/rIK6ikmr0g4Coiic
7dr7y7CodId1wrkQDUfe+d+LM4e+Q4uOgpwrSvl3SNu+eAXkpP1sJI+vVVlKdIbIBhUXvvs6GAeC
zcqWx7G3Zd76DcUJ5iLI7bjZidGgPbhXmJMK37F+GPXKggOLdWi0AIfNwOj/JZHdb2CbhtH6DRmr
E91fuOkn9K1qen0EUg0qwHIMRPIyrMPmxSHI6twMYw0ozaDIUdkoMfum0/dhNA9VMpwnKiFeWDfe
kL+S/+GywFgwWVbn3j/Xns2Je3Ncsc1K03IaFcbt/W84diwW0azawKeeXNXRKqIbXlzBE4vhaqmz
PVGmmnyL4m8SSGeuaqwV+HMMmbFKP1tpKZAxR7LbHBQRAIh2cSk45VMw8Oal8QaQyUGqiTbMqeBA
e8n4ObEecP7wM/qs9zdJLzaYoigZ3DN97KnA/wRgRrmmWJhpLwUQG229YS+4Zw/3uysMIhXbYQZT
I2Yqjw4XpK6/Jy4i3MAvKCV/RrzW2/+YJY19GacbQMvL/fx+TPE8hgJz6EFVFvoBsLfOwsu7Cinl
wPjrYuY+mbvB9sX891Rg1EKL4X4xNwp/eKuES/ZiwWaSUT+D5EgW8QLg6HLFm4yp4zW6nPkrGeir
7pp11K5u9U7kdwsTfMjhCaiGVRramPr9lP28/nDLu5RERbiFC7NqwEboa9ghAi7xnHvkhKqWORgu
8M24VbWR5tFYKaj3ds+rqTH56952BM4v64eZSR1ZrHA8+ff7OlA8FJLogq/dcsQuyKL6ORPhlv8t
uIGava2EGT6WSUud8bbCPC5Bt9/+M4kzEt8Jai7b/b5joR0bKdVwq+uRs2j9+DVPa827q10lo3ei
GpO7ScHPoMuMk7t/QpY1uTm6yLD9GS4yD63yyreGBumOR7P3nTeW9h1/La9kiSZk3NwFpzaBPPfR
LDIVfnUpSKLU96q1F+Gd+HNAOevb3kcvvvKMjMV4Ua1isrVcXb0g9NcOVyyNqT9cvE9GUCRxglRk
FmELL7JMD8VFcAK0RGINicr2oLqXP3yOsAgcO6Kkq7EuPP8iSR+EDyQIVhmg4kCKtjLcON4hnV52
Tp0xl4bgz7tvS4+sP8/lMO8VBAW/nrePqf2uTfBNpG5FwmeqhQ+Xsuxq2DlYSdTz/pRGoNCy0L+q
Sz+YLlJv/oEXQLrNLnJClDY1+hOmFOTKK30UElgo3MsbNysb/HYlvwPRxjfLwUz1DBIoD7y1M+Yj
UM39uwV0zKtgIOECPK/DazpTPnbLJKVqGE3kpjFUoenw2Dpi/qbVG8zuOdZOZyGlRwtPpY6W35fc
ojITNQ93prkF8UV7aww9ZgrTOfRVuPAhIndVSVs7LekuCFW4G63fhVIdKqEQwhVVzJcmAIc9J0jp
bKuK5/KSIuP4RtJPv80yJExYEDiQLtiQZZlkxdzGYhM/2FajhiQ/etpLpS/LJfDE+eVVRXsogaIK
9wIAzx7v9giRPh02Z1z8O8HSZZT2HfN6ETM+Y3GMf7+9hoWM8vfQMeHbeLnX1usGy8TGjDDB02W0
MNcQH821gezO+OCSmM43f7hKDtdTKvqv7VyzERcR4GG2AqvJCRZf9LagSXI5HLBixjuMhs3SB7K3
V5OjVFkHtZoHBdbAbh26z5+n85EKBE/9PzEwP50JnVGVuYCJJXREERJYmAjhxaBgnbvNk2gYERpu
F2usHY8yBaXnqzZxETZCQMxMxi/gM4h+eOQomkgkg2Q+NGK5DwW9JWCDAAWJEBABg4NzNJyg3mSC
+Nu1/BIoEnrzoqo/BHekSIi0waes3i0qmlz9ZDHpb4W30R2tQ99OwojHR2eyRLCcTj/eWHwRn2nY
AOMhru0nRPq7+fB8zpdiYSemBucpcpDvbCDmCBC/se+Am0lGWNP/4Ky7BZ+Pd1+3WAVDBuGp8gYM
vhWFgQZCZGj9wGe0O9YTM2Z2JK0Nmf8A8GmwtAJY3IfE85nL8il3REExUhaKBviSEBxUvCnfqGWT
Vjt/uCv+gjOUdxAH95Ry/dGtgGgmhZKK3+OAE3eo5MPu5DkxkX5/rCDk7B8412Lvdqhryc3wsQjl
KpJX2Ub3SKrlhDTW4CY+7g1KzxMaH7Vw55tdJCwxakrpjuinQg3oGbWrBJrMAycJFFF4IJA5Z45L
xlNBYFJPzgCWmI6ymiO/y28CiMeGFd4XFjrZy7cH21i9Y+S7iKFmhCqv5llN/CpXWIBvTyOFm4p/
2fRt83lkswBokGazgwK3ZEWn+GoM6ipZ9zrb5ChXwHP6Cif7fdmQhjODTMFYJ4mhLHIwubn3wPmS
CdM/AD6gy/I10qKgleT/msmjmpu96KNmkMimHY5u6xm4HNXqTXRdGYY4EKi1Ui6XdnRYNLg+oiTS
A3kPfwVfbTjmUx+mT9A+3mLWoYPw8dYbBjOBt9DvbNcudSrjWYfwZZt22DLGJUVYySXmoO3iRa7G
6QsZa+t68fRB0JAwaFhRXw/eCS1w2bhLTgEvrGbhdXL/E5oD8WkyIpBbMNjUlRhD1SFdBzjaCxt9
D8T5B5jpio7gTQ4CXkxqs3U4RrOGLN1iL4SwuEgF7p07/fxnt2qTVnldPsenhD4AoAQVjfdLsqKB
SRImBEmiJSSLoM5MUyu3vBQmlAT3qlS/XyIm+Y5sLOichiIw8mDj57FMzvHyZ1XrspL2CTOqJ3m9
MOf0CnKiR6rIFfU8+4OSgz/AJWLSQ5BsLWYGYCn2b5N/xLe1dwBNVam5BQVAhS9omj7V3nwhuQvS
VkfRLua5J++e4Be3Yv7211I1dPTRNN6rgZyj6fM1kFAqx6RGLuFczFcC5qagnCTZBk+gEs1HmYpi
n/kUhPx92anxwoMTFp8R6KFQNDVPopR26r+DVl02G9zmwZqhZ5+YYiKq9BPqfxPXc/Zt/WxYnMxX
IrA/mTjn8wI2AioEbY5uzntrKRlJFezWAStKEiLlShkBjuwJ2NBR7D+7JTkeyGhAPn4cm5bTlp5K
TRE1CY0T1T+IRc+MMgeIjuRq24nzTuhd1AZXFCxR/sMIGBUwXJGAiSh9hIPHIJAOd8txC6JhnICH
cqu9vOEziWxVadYOKmwVZxSqGQMbDL8/Ers/siQwbjLnlp4E2U8EWOEJsQ0BRMsGCKJXbOgFC4wX
g6Uk605FFDMZAqK0yJtXE81N+iCKeM9SHtaRX1x8sNlrCA/Ybg1uTWgE6ItZIbjnubauKtail0V9
J1SrIW4ItWwF38d8SnL25i2ICxim8Dn4QD6O6fgha3hnUwcncLd0Ai/5uYl4dQG+opBvdpI2Doqw
VznTFTjHX8HjytL2zGBf+/1OR9MoaRRuBeC5949O9tuHwpQaDYzj0PHbaUt8z+Q167NfuE0q+9gD
Nz2R4xYjWFD4zErv5hPGEnGlmZCr2OnrPTTytFaFgtlqugIpsaUDc92CxAWxXui5Rd+KzPmMXcCP
WoWgm8OcD/v0tLUD4iujor69dzQliWWW4miT3RwoPJBnOvFczzpx7As+v77yTU+3O7iEWD5KjTLJ
Vzqsly/ImXT89O4Wv+46FYJwE6G3X2VD6VoCSLUXp43nCy4Pn9Qy/Ssfs9ro/iAd38iXELjuaY6+
+q4F2Uk2Ipv8xKBTHDGL5nvvTXckuLokKXKzehaqbd9DIEfFJgo4enTvP17T7PLZbEAqx3sILz/4
O4w64GqsJ4yrgOzhqRq0Js9dq3hP7wpNbRi/8QnRGtbnLH17z8772NHnO3FH0ED9ra+/ziOP2IVP
LZOJ/uTJVWvnbTMxBJ6C7EMnHE7LuJccLp1b4FOEjnKA0GfAobACZxuQKhg+rLpPaX2og87resRO
HC4tIyqr3cT/Dbd4f5v0uBICBviFtwxWoAW4VuQmMHmCWzJW97/JrVLNA+roEFFO5NIJ0hnyxfxS
aCuIZrgsqXUKdrj6quRyFlvco/9clyE+jnmQmaiV1sbNyfkD5wf/SFVr9jrESV+Z9RvbAsG+CKa6
XdWEXm1s5yxHnem4uyT4QcdhQoeymxgI4wQ20hsNmFkeZ9ObwspxakhwzPImgdNyl6kolF/p3t/j
tXECLIsCyr3KaTHetObjdCDEtFouo5fBxCFU9QD356coTGqSOTAqAkgIve0nhOiQXNbPT+5aEJ1Y
NOcP+tZN4hSjvpiI4QAsGJW6XGNYLT42VaXWIQhQONjkESy66dNoVN1f5sLQXZa6h+53J748abK/
UGj44dXfsVzYtkPk61c2LNTZPST4PMOr5lgvISxBnhEWnhWw+HGJztI7ZoukJde/ecysy7JUXEmg
keUpuEDDDdogXHw8W+p506K5Knu0DqnW5aie90suzU3RnbVqeaUvrE4woUoQI/wEUoWM9L9hG3Q9
x7rI3oXalzai0ocJojf6Pqo4XWhlKQNimQMOyREzmEN4XkCH6DrDPoCUDyF1JMLh5sCHw13uGlQ/
/U4GM78gJvGmtCRi/y6qItWnpVAIw8qL1Pejqip2RsUyGZQ2duhATi+8K71Y/XF083Nk90xdhgAN
hZ7yQ9WjVkdODZElkRo/DRV2jDM9ilsO6w7b+vMt9FKfxxZV4TAnBy6qBuTNp4m9WnHwZ4rL05hO
yOvbUUNMui6tO+CJzRFRliq0dInA3/dcOGQWSUIgEwG3c/MfsbWtephwLwqdB7nvfJ7vYZEOvNsr
4o+jrPOhtrMAunn4RAguVPIzEIpesjj0Z7v2iQeOw5WdUUmmvjigQW/Ypn3sYJDEaQPes35VwNYO
q/iQdm5UG9lfqSho+Bw0pob7Z7pLUsvTNPbzudJdtLuIrSPQVejReq/EcGCKIbed+Bex1n03uwb+
kKRNXPpovDAioq3OE8TMqtKylw/5yxxUlHBL5smtqhf96hw09XjeatQA3l/pgBJVGMaDQMv7l2Qq
jXnRwXab/9bekkRz4nDjQFgN6gG0+HtIopqJbh/vWHdnGr1fabyuDossYSDmJbcIzBkCQp7dnlSW
cQUWN9X8pG7LgKIAgyp1Ex2IBT1TUeZCGoKTB/YNYFQSmE7EkmxuXhzpwlR/rxFq80QMFo5+GRnk
SKL7NLWwNJ0Q9Xcvuz5SpJmAfw2t5oNVtbo6JDs7iX0/jQehqhue001oKkQMwoG51gKFSqaxDjrO
S+Rdw5ZrVb3lY4dNlDW4xpQOoZml2W4JVVJdpHkfjBvER291QKnhaKU6k83O20xLyL5x5/+NNCBa
ZFRq01zxYPyiWP2bLM7VhHqBGeB8aCb78G7FWXkxJwq0xUbNl3G2V/euBwpShxBFAkwPpgy1YYJg
ZeagA/UIHphe9coBEmxuE4onNFLxewgaseM6LQBfHY0YYVoTWgahelPCTh9TM453apUbCvO8UdOL
NU+Y69hfDMJCO22KfBCaR17CKuNXB+3O88xk9CpdEpVHoCL7wraeoELqTTk8Ufq9vcInMDLAvQxs
K4HHdEKgtmrTcfHhCorXbUYT372oaFva8TcE6EOXVO52Uxt9JY7E5PmB7z41mz/iMyS4upyE3ed3
9BCKOvFfyj5DX8fvomilMIiPdj0mq9lHlPHH9C+7dlnVCLJQDOW9a7gQGuS52AUGmBuiRsfxUujL
OW84mX2lSzT9499YQ4/vVrGXqYdTFZgi8JHVKwh56xkRPLH2WdqP3P5I5kINvdGyJpjej8H3Xxnh
sGHVMnXvqBulU87+3gx0PaW0wHm2V49UpwBR+fxEr0JaahLhWzAxTU78E1nK8A29FR7hUeXI9dRB
zXvMGgaxGE5DD3/0ZWB9zqCASKyzrpys+tqjZr5Zfwl6vbmgwKw4APxgX3uyOL0CBI7IMopP3AbR
ruv58bEPPjvBGrtt7DM9zznFy2xNEjxX7eXKBnLwhRPUojriPFcjhzYP3mz44BOzcXaTKDP9iVSJ
kfaMtOGJ5V0c09312v8fs2fiNLz3PbMM5fhsSio1i2sN/GOdAjfr+eKLEZdi4w6gqaSJMDu7J+Wu
cvm0rjcDHk/ShmoA6w5BrD7uO5sLTnMPCpSw8w0vQM1xpBe0vrLN9GFUER3JEFxQdCiBf90yvt0/
0kerYsvhdbgQ0cZnF0++XyYPMC+f0wXoD1bsO4kkimm9JVK0lr58GPTakJ2vPWfyb6bJxni52fyS
cQPw4wKvjc6jXTJYRuXk7KNnK6JAzXw5n/7BuZ+a8M30Nwml15uZb1yJYtC3Ieh5sVZhcZzvigHq
o6umQnVPrtCvqo2gTtu6va9P08y6enGGCgZ2+S/3IZ0jrU1yBIvHyul06TYLJdGqew5eFjxxJpC5
WQ5tr2a6GuGivbj8UkrNp2x/fN/iM1VAHDAM79YDtfpoZxk5Xd0q76RvtU6Q/52W0c5b4TuO8CG6
7HGbiKHhqgfLRFcu531enIOoy88X1h8pNKGm+cKLmDISziOyDVff3QiP40JY+rEVWQ83vrrXjQyj
BLPlheXbgNmEiQ/klhCxEOSYxuo+adzz69jtlQeqG9JGKCo7rsTeTPO7MIJQt+zJcpRAm9miOQiM
0C0LMlhGBKxEekx5C5bVxjTTPE2LQu9pNINkTl7kYmo1bbIeL0+zsTAbghMVzlIQF2IaSbo+c7dc
dXD+tA7Uap0Snxrvsz0ce6yhgtmzAVInL8ewn3tAMaDw+cFicuxQoU5SNeOOYBqgqJRcxXI/9irj
yMMvfvw9LrvO+Uv/OkmiP0mOPLpl00HZQS5VFYJeDynMxnaeGjsTY6Pk2soO/fOo8U7sdrphmmp5
PbHblf3xDjXW4sevGVy70KmOIksb1TBpNvBDHYiFha1nESERe4QZXkNaS7fq75MIH19iiFM4AOqf
vD/LqP+d8wVNWqX+LUMW6OytYLSIh1yAM+mQR1GuPs5hi+SMlI7zwcpSmnd03TSW6AMdkUu6x9tH
nN5CLypxXzyMZ+6eChInfJmv7XKzV/4Ep64TbVSiZGiDW80fxVGfsDlt44cCN+RzqWwQU2VGAPAw
Ha4UG18spcqA/VqOfvpTyKvT7+PA/Sh4wgr0e+HMiK21oZj5rG/vP0qAEjvCKlA2OYehkV8jdwQ8
FjnmixGuI+fiMS6AY3T1rtrONiWbYZbLY7KMd/vUS9xQUbNdPYnZ6Kal6cAVbcu/jQvu+seLY3Cn
8QoazyB47aePk/rk9hxKWXlQaYoUqXeO2zhH6BM8CbctMXePWPATJObadJrx2+49p4cplIU7QhVd
/o2Smtayp4e6hpkuPSEKYS3GXeJYNIvImGIaEYhemhLezCk8F2DNrdDX5NphOxVNyxYvBHy2Ta0w
HD8SLpxf4by99VR2TNyUAc1U9LwRgJPVa3MU4Eoss7ThlSudpFTMgbPXXTDHImuuMvpk3swKnCD8
nhCq+RgTVZ3NeiJ+LatKc2QWb/KLRlf8ZoR341dB2CQtqevDcetrjl2g1Z+/wqUdegTD1L1YbEFk
5LqCBPJT/LrUMdbV9XQBGNm/jYBc2IIXnUYBqvD5U347W0Je4nMhY59zk2OuFedDVnGzwEGeKBYw
hbQ3JE2sY7WawWL5Pejshw1ncb7jrtdQfP4OUTDhzhYoXrgeCQjha6B4uLrGHN6NF1UmEVn4HjxR
qj2vL+IvS+VGMWqju3XlO0SIVc3jBLnIUq93ozdSMktQtCM2bKcqWTTOUESVcdj6hA6gugXAEj+b
EIo+RoSM2XBL8IDnyFTNQ+/fl0Mi+ceinvGxB9bH5Ii3WaxDDLTZp6Hx2+hFFXm7Dt1Gliw4Iox1
H7s0KdbrvLkMFuig0UYNhS8BvH6SsFg6N/VYQgYiyOZF2zzbYacqWyxg0+UW9DFU8LumBNcRNXOF
NYiVQFIbW+tQsUF9+6Yj6gldgycvcct34lQY/df7X8wB4B/Tp/WsxIZtfm4N26U7deR9IIGpzFcL
veYeWqbCfAuKsQ31xRn7sjrgfhOCNen6FT5NklVqEwCoT+VgGZgu3KaQqz6qGebl49AI4LpjRA3G
4ctvyjuhV12BBETSetak7FJPbFDViiXU9UDS5YF+ASWPMxVusFZkd34W00FA3C7++hdheNie6h/r
j7tS14y5uRXSA6lsR+K26WVwUKjOdgCM09t0KZWIhjQ+kDzcOp6elnxIgY/o+yCA+NznACu9OXpn
dt4orPMa0JNcjanBDOT5z+iGA8Y79cZ4LQ0yWNZ9bIwq0mGo2224AomXao/s0paxXT/gCg0GtQ23
z32d+guJIoCl6Nmi2l3dudrirgEZjhyF/JAROyvG6JiSJaE4CWjH2V5PLq+Jj8WmTuA9TPL15kRI
r8IO+7q7uhsXIvbECU+eYwxhZRifp+KTCQgIGb0yttiWqIwZ+GtWtovjaipx6HDd18jac8UXw2x0
8jOLRUPYtncXIPXM5HoO5J1XyoWDgwt1kA1xOU3Dj8QFugzZBnhUNayMTCbu8AG6Fg88cBWGmEkF
kYodTLttA162+VjgCa/ILt+02jKEAECvQ8sA0HP9f3kmTbAavncG/6Ygf6f3kCrzfZxyfdTRkFT/
u3UVFep3uDAXR12QFksmY9n5JGBfcH8/34fV00ZBmeOOaJ2V6x5AImZU/xoyTyf8N8YxQs/qwVRn
a2PnIY93D3T7D4jS7NJEZiPJTqB3dBLQd/r5CR9p6B2tgPWdRHGh/bpUlXkeLEwwxEaxmxK/emXq
HEVjvPuBMNThDHemFapvZLnU2G244Q2I+7r8anDtr8PEidb/wTnQ+G5tDuBDuknf43wpJyocjxA/
IwBVxkcO98hhnXLO/Wgx82N27xUnwQ98ZJjCp06RFK55UYk4YWDrQnyePpT3gFy4tTswg1Ysm3yr
tyFie9pBrFICyt7OlPLVv6uFUqaaTEVCZ1hiq5Ypfxo857IfOIm4tssB65USCv1JDhY6JYkzVvJo
HQ4G+at06wzzKmXnQ0ubTiDCHm7QdfWRdfxnw2jeG/eEMbkZcRGoIDFI384YmN16NZYKLQD+w0DA
BjFpsnNfX7Nto9o10J1Uar3vOF5OWhG/vJLDeBIS8w0+43EBDBk5uHphv78abcvkuxwG2sEbZU18
DhHwz86vKAlKJgo6tPlMqfWcceFIECGngv1h5w0jKkiPREeFIzbALujPwIDY3Qh9A4HHqMydYIEN
ca5Z+r+6kWbx3hw5KEgXDhyOCzOggEqAwVzf4E1GOztMID9ki43GInbcd8t+pYNXe13tkW3g9kL7
ZZoisCiWWyOOU0xttaUHwcq6x3J0/Ibc9O3RM7q4pYv+uIP6SCXn89MX9mBSq6NY0+Gh/nlokXxG
EUqDu6j708XT6q6h80aJyOrzd7IcufINu7tMhEOfcxVPFJ3H+lji/hvWjoDzdxpMnkgTYtVDeKB2
Xc+FRut23/TrrEIEoCFcbXZthjyaU2YNnL+kYOf7Lj8j1B6QANF0aUD//BvkL/Mv+KvdtNdzzFPX
A87j6K7SJ5ZAvQAnIO+6jqWxgA8vlJOtMGiF7yfb8Ewycm3cc4h1kQZuBsNVfAbv0COquHLuH6rJ
i+Gq9FnicA4iH+oeUGrRmA5M2VvE8qBQJNGjXe9H1j559FR3ntGtT5kmfADEZTkcRvARNa4OlbTU
bemQEHgDG3H+S/g/A/T9JkS0romKp8soAgKex/bmv2DcBXiI5YljOcDQawvDa1gAht6WduzXfMz1
LYolVt17qV90TbQOSF3iRgP+aEV1/wNf7nWeC7Ed8/1e8Lit35qtMpGreHVX9Sxfr2msKnGeR7WV
orgEr8AlnbL5AXuf3D165OHGFZj1k7J6cPGyzjHq5168mv7dbLmK4onERGQepsJcS/DblWLp/cU3
E+wRM42+MpOdQuM1WoxmTq9kYiN1sYtUU5oguEyhXv2Sk81+agbFDoThIZgrEtK68S16ll3WpzJz
ASv4zbSfhrphKlRZ88gLydwnTh0+NU8Ol1gCyrgdz8YJsvIjMii/U5uZ3s2fQIbuTcAlrAdA1tWD
o4L++HFZXXZconesXN0WIagQtzE8FVxWdd1athR3woMvB/zNbFcZIJBlNz3R8XZJrGmxLvNNydXY
Byr0z89ZdV9+GvWduUDv/L/PqH57VR32pwv3hUx0QqOaeHP+W21tEeGlibaXMfUs8BUyV/rH9ULJ
hMXhXMuabExxvDR8xlf1p314AxW5GhUfW+4jdZs3Bb3OM+Ue6h/3DXB9qpzRRJbB8zkG5toKiOvu
ZSBX//inOp/N6qqSn6eRmC9YX2IpSCDbmvCWeAWBoKZkzKoqRu73uJ+aPL/LYREmMZXvNsADBJ4/
QjXbWRBNrofAE1sV+3+AnGyH6LdaGg9T3mxujQTd2S9G6iTxe8ZjmkzUoQ0xpCHrsnMQG5/bzQ0w
Kt0N/oZE6vFtYQDnoOIJZcaGQPjT/ds2L15jj8CdgC6Zz1kjKky9ZAjpJbPxqs7lH3tYxTN2pWrT
en4C1wShaTCNX8br0La9GH8UmFjMszGkpWMncexQoZLZTqRWAoOcl4Q8hoSWgRD1zoJ9FwRbSgGT
ZaKTX3zu35La11UEn47Gyzj/ZuzaURo5aYqbFW74xaTPwMxUPSfGruGxPTWhsrS3GrWwrlghga46
ZyFoOqoYoxus0rXMxHkgXP+5RXVWzhG8g8ciCrrkAUlfhHn89p7B7aj7/lTPDcAeuVCGov/7aonv
pWX2hATa6D57RqEunsT1QsBqVhY3cszungbuJlMivYqj5/jklq2NO8EPYcj60lh5PQQG2tJaqCN8
omKNZk8jDiNiy8hS+vmZlPKIH9cI7pIsfYQvh5AMknfXOJrhsW14LSIdOdR8RwXZZ3NVi/I93Dy6
W96d9vuDJEkFrPdIdQiV4rNSyNXlBZ7d32KnBXdUJKuZ7MbrgmZVeCZHtk2aaJ0EMfctNeUX1YSd
Xxwl0oX85HdxuuqCZND9bnFbsvMgCapP3NWy/rtp6UZ/2Q1oR7pzyyUkCZcDjtfw/9ft2UovggZe
obqiZmlAjkq3kU2s3wiJgtduWDQeVh80aK9SfbMX1vMUwfQkT8wfhT0IAF7KoVMe2YweA+CRiKzh
HuoX7fIFiWhk/y+aQkhphZlwOnMa+1KLLTExCewt7oiKiaXhuoRfaO6ma/U5p9qvKXh/2KM26jh6
PlnDIS0oFZs4c+k+RmegVr2SbwLifXYJuosbRRcpyZl+gb9t0WAZKRmYZXXRBFOwGA4NiF3shrgO
PRt1ibZLr8tZW9Zfs0zg3qtSCkMtris4xR9wejDCKpNKVf4hfq2Z3NKSTYGT8t40+AUaim5A7OxQ
KQcCbIo3OpN5Xq7DmBNnh2CFsAc9mTkP+mmWHiSqQO7P2nPpNBWdS6lMRRBI6xaFk949TPxSRPwI
O8dkGxMA6Yd6dJlLBgrRhoGxeDOJSv2xbnHfVMfRUVilUxXOrjRmzv7st8o2xmyltVJaCXlBIg3r
avVJDyj84gn5LfAeLNY86Fe8Bb7I/pSRghbEJ+eXQ9cWHO+uDx17Ty7Zbk1UHBSGEgW0Y42A43D5
REh0aGTLslt1XhAYMogyb1g9WldpgR6mhYSkqKwrq4EIVWIPjRXEVZ0Bcw2Z3Sx6nl+Nc4HCcxsM
QPZqmFzoPvd9YXVxu8FSjgZd1zSXnvAK6zUlCL0ZU4vT7cIWMe8MbEHoIsCFMMCYhDDHkFX9XNA8
oH6XtRhosnOIX9DVJhhAML7U9NTlRoluP+6cxklAXiPtMVTudp7o573NGkV5TYau7h4rzH8wsbzm
YcezMqfbpcLSEwtO0Kz2QKEQk8vln1Ozk7CVmYQHklca0sLO/WFVIhvEi0BABwEgkKvZdmxWL+9Q
BlpQnRj8SqoNB2zvF737W5rLfu46aRNtTrvsi6JEVh3czRJ1Zb+9wRklJnNQM4Czc2ArNK0UI7AX
+BMIw/SJSD80Mg6K8LNOqWb/jeTxn+fqhAL5tp6EUe3i5dsXrqouc2gzQw7mV3yGY5P/2yXOUbai
6ubyi2o6c4g3TNY5HLyDgS0ozBUuGyc5qINmR7f68fp/e1RHUhTVQ1+QrpBs4qdgXdjBIlpHbB4v
bt4VB5d/OOokJFGwOAeSmMojG+2vG8xhoLu23pnGmDOEpiYPaSS+FlaKgorfpmgQsQp8yZyOzhAO
8JFXoQm1dGMLIn0SjFVWjfm9nShFqagVbX4AbqE5MRfgSsoOK1fBmRV72Adpx7aMLlxixd0ndmkT
0U88Yp7dDIsycfbLdnoNu2fcYqmaSctXOQk+lJQ9uY211114apIdjRpYEvyO99A8GRrs9ThAsfp4
XdsL1ZES9FUE2wx/6d3j9gA+WdKSqweJsVz7RD/uhLk9xR6n/sc3a7sYhV0757jd2oCAhUSESNjm
KiY6LxmSOUYTgjB3i5pwxBn0bVSP2A0tP5uLtgdiyE5W2+zkdFuEdyqqE3Bm+ReGFZx+yFwruyRw
F2c2w4QTsoXwnZ5YbcaTkvrMZScDyJ5rJJS5ABbgGUNevN6QfnCM0XngsJkuhynDbBdZfWiS2oL4
pwUGJ46VPrvk98i81mSVanr5BPVf2WYbT220szClIuHxBZ9rV+kIpIn2KcxGsMycK0UeZo35dTBo
R3+Qyqkpn2Ku3By3XE65L1pr2jaMMyOHLrntNfHOgSA4LIC2N/s2V3NBnjaraBj3yDCbUwa7A7TM
UgINBcAKFdevpVIEBB155P3Rce6wJs9YpMr1qdBOND9Jam3P6JGc/c9FU49RLSCHwbwlbe3osaQe
8CIY7XpH8npnrlWr3VCVd2eCgdcMSHfnSAozXOB5ycP7Uk7KMQySneEabIS4qqmZpNOmcvA0aXn6
N1+UPVhd/dbyiOww7UL4fWGtxaIU2CKSrdjbpe8Uo9fNkbDBSDHQh4V85ZtxNeDc30HyLnSVA1nJ
zCc/jLAtCLd/W5m0tUp/ec6qjpE17zjrf2n/qM+O+RzyXHkhRlPDyX12Jr/O3jPndGHkNRzfSvhe
mMT9lWItAlEOqj4fOwXsid48Yhs1V8OdguR4ag0XS7MNOUrIGu8yvExmrcSbLtAzxOnZC1dylQKX
icnlhJwgaCwAtcRfY3NQfR/uf9X+M9v+leFHwdKFILsc/GlSuqzPx8IEwPLiGRAdMpAX1CYY7Xpo
kPmWiWSF2UUzQPDU3tr9+I7jBxsoezq0IDrYPbFYaushIV1COMVWu/OdQhvXusZqU0RBAetQxAuf
5DXH6kaN2QvD50sKQLgBB+MyyHjJJzVhV1gqjMXcFomQdKArqTtpDdP/g8OQlDYpYhn23ug7ab/x
3p0LnOZhXavrz86irnk3g81GNew3ZLsn/2FQSdd0I/WTEf/navaB/GXZ9y8S7x7yxes7brOFZ+oh
vpZ7lTrkspTeYzjzkco1zYS05LCuSwSau6f2i+PHd5kk290unlfoxH+Ub+1rnmlPnuGplR6cUVA9
N8GkAldI+UUKMTXbAk1GPMI/Zx8LzmQfwbqQrjmb7v6KfN3WU7lrj8aCKJd1KRunptx0N4Q1+YqS
TNJe0DgIWAjw9RDu7iUgJiayZG4mlefDrY7pPww69owDQRnw6ODBp/3fvtguTnMosmMv91pyXkPl
9lHiPEm3JL0Y0nHBs9IJdbNXqXnetGRivnNF9iaYS+LCXn3/dBQ/nx3HfPahg4tS8luXvaoLXhQD
BwXqTUFzARWzBwNWERukxO5sqbcveQjJmCTTW3ZgvM7c4b7E/9m8qCpsqSG4FsjOCZL5dWjTrUhf
x24NrFSwyA9NvlOTo38IJraEugq8nH94JxrfhGB9fA6Ejprky2gLvh6aKaxhpLhNmTu4BDoClsjt
a44ntbOHngO/35EHpOmDAEnEyNQByEO1o5QVdlcKUeAtg15yNMZPe833JMg5uE4BGHMuzQfEAZYu
b7U7/v7I7EGc0b/KfuBrv9UTfaQCfPycw6co5anXUvMEHwl6sgxjUaN/Jd2of3Glzg8Wm47t47Hh
IW0jO8TC5t+Lmmoi77S2xCYozhJ9T8Xy+cQW+qAOMYaaZGVaGOc8KF2tevc3ACS2ffwzKc0tQHmP
iSDwlA9ALnr9jdYCyqneWJ/OdORI5BSM5Et9xG6Nqkh3AHLl4HzLd/vnYIuaNFzv7soN/uOpBg2+
3x8YH9cvOS/NDFZIO8/4qP24o5mnAzY2WGTsx4dV3Qd4QQ3LrM2FLLUwXiXMbtm8pD5YXB7kD4mE
OKBSkwWTr38IO2ybLzKvGxS1FAiJIR2DZzgSvcggx5uYhPN0U23NcKZctqWRpWGmwxLjUApopnfN
2xHHvxe4hbmRVCY6BaNhkLI+kj1MgjkYBOmgY/UBb7zIkr25ZqbfTSenmQjSf00UgJsaYdeGOad1
ZWCR26V7L+dxL6IcUjfZLV+bv1glL3yeuK4E5TyxUhvDlr2GbRfbMcitMsrr1IwWdW/UFzwIE+dT
90i2DnWMZvx6x9W4pa2ohVJNrofGZHwdHkoHY43X8UJRYj2CTDlXFt/5YrLWDkwx7LDg9oWTwH7N
rPre42AOLRcY2pQnLQ7z9dPi6Q7I+BiEkgW8BTqRTILTvkp6Bfxv8mZqRi20OpQRqcdzKUdjUK7p
P6sZB0e4oOX1YF1ncXrnJ4Pf2pP4SHPXeACVQ0OgVbcrv6p8rR9gd/h3+uaZExceApnrzIyXECW7
Se1j98WEkzwWwUBPZOkTWgRaUkUe9rbKdGY27HaSK7lUkuBibI2fzQ2qOMS/+QXUIPs+Dl8fAJ+0
p1kpttQXlXmqdhxvDkq+L5RYkV94Hh+9SC3qMjMVA27gzqUaxTal0Wjaaynhf6bwQGnK6sUYbRCl
H7ujQr5M3ZDOskvx3jXR1XF4pg3oL4YRH1DeTZUeXroJokqIW7/4kjS8L669ha0EsVw21SPw9iNY
SAJRVKww6rHZgZ4hU/8LRaNO98gHhw8fSgJjukWs1Nso3g43fNvoByszIIgm57jksfrv39TE23WU
ZKVh7Q5Z55mXhkXVCf5RbQ0rZENAFZODywyifwlVVJ5qYShrpiXdX01T2NI6aDYHEBqMGMqwM7Av
De6jtakV4VIhRVxnF7OYQ2kSpjX5ZUtdBTkJ0gSnezoQ8zSN8VZSs/tlXOe+kMJ4mRhCM3sXpajJ
eszx/oWpM+PQC0jMDIXU4k/cavWseOm147BuB83KdTLgtkJuDXIMZ6rREl8UAR9lw7A8Ed12WTCf
bJdv+kMPd8Gv2dEDnXqrWYSosMxrXT+KYgl1eVIiDPl/63v3xSU78P0t7lhLBmdgWg2jA4mRky2y
4uaJe/GSaLejxnXbkG5DLajByV5vLDoLAgRSl2iXU1milZTzcZ94Rwuohz6Oy/fOBdd2DmgUK68L
6qDV6/7swIEvz+tw8QNPlkukCOXStmeLcAYti3UUW250W8ErziU/HPOHGIn2SZr5e++Ad0sff9oL
eqoMuj1vQLC+mVYlPVEEFZjt72vJy6/6opvWwSlFmlzimELU1On8vQHjpN3SQztoNZAHkcHjC1YN
7BRfGKPHJ40PisogOIrWMOjaq81vKdSDUmf0P/fgOXhUKrZxHtHXPHEmtLGyMQSJF0rbxS+J4yDm
VHZoyH8LwO73Msao2GcqqMVDi4tPVCa0AsYlpD9Ami+2hUOcfrnD6mVqGkWEqVTe/DsmelDDHHfE
y0nt9wWsV8GIoGsLc3o7hJ+R155DL6CQTeOMNBU4+YYTm3GYGDpS2jQ+xTs4CBVK1dPmI+yBair7
X7MJInwxkRMlz4BlIe27sdB4mKrcDHGZR0iQNF7OaTNV78B0e7DYha7bmLQl2Jc+V4UFuNHUogp0
JRivF0CeTCN32hMYmfHMNH5hPJZ54KRLjRuHd5CqVAAGF7GHb5xHKE8Mh5uNlyqyWrkWt2t1Y62E
alSBR5Wt+TzctQw7BRtXTaTu7OJ8Xi54E9v9UxOA7ib/P7B0asbkPeYDQxyCiSyvvuoWhnQu1od+
UCXOB53Gqv4Q9uErnUJqOubnP+IXekA9aMVKgZ7BAqiEIiw7fchtg9W5oi03VXpGUHlsdU0WvKKt
2HWj8qg3sm50UvP9DaKi87Yf2+WwdUmW+50IsSFfIKV5UhzqfxUCZFlZV8Zn/i/NV2/kMxDyHfHu
oC2VawlftcNp0QTpW3ZYWhyILKv8zxJIHw2k7vrNl5Ie3mcQV+aTgUt65yqaeIpldZZzHrq7KfRw
2BP0XRwAAcHP7jvzIYrJpkaH3xPZDUseoJ5W+75CP1btqrpLMReCjYxs2FdNn1CWBNyxhf7pVsZf
j0C9qI0sICOGDuKtDLdJmPUH29vFyUc7Kn+WLMTAR3S1EdU6gcrnwp04Vjs1zL8dfyxlqYz4G4aK
+jmXQOzJCg4dP8NyipRS6/2Qtomi99AjGTCs55BICQH3tNmSC/4UASWw0OXBfgs3lWjNyeC/J5Kg
3LmBDfdlnG0wUIeNSa+89vXnHUR39qoUsm9Vn/DJB+ZKqrPX1u3+yl7RNDFhP4dtEnGCSpphb15D
E5kPFCD60Lgg8usQ2SqxtBY51Mh9Dsnwqdxnsz12xy8ZPPyO3tC+haanA9tA1H0WlAU937IEBWpx
skZWoKLiOtE8zx7l5nIfwpC0xy6u8CXrw2/GXaeWy1V6bVHFH3uz/ExQHcjF0XE0POeQpermcGxa
YxNCz2TCZ284OqnbZ8Ul7iyYtOQHwDqB5v8dtPH0JqSSF2gTYZWQUgLTbpT0RSUcfTp+GRiPkPbb
N+Sw99Qk6kWNz+T9oU4eVJiaCRUUvk/LKqkxBeTuBKp8Hb6n+69LJ+9vEiT42DITYh6efxX+mmB+
l5fIBPBu6F6Rk4kUIT7DGwQHu6Cu8wj3LhUt1pNsjNmKT6gTEGF9SuAF4NgCuvLK84x8B3QT82w7
x38nr9RUr+QR9oOu28CwAVKhCXAt619y1wfm9vRITe0/SOLSuOhBRWXQjQ0i1UuCjJfMI9WWl+r7
Ksy+bG2fvlXtF8J180QnqRWP8b/3BfyLHmFNkB1L7n+KUrgiYcHW62NDhwFdLgGWeq8s9/ncrzl2
p646MYlsPUlw1rBl4cP0PB1gyfJKYZnzPkNioxPB0FKQOpiLxyR0aPfVm+rLshppHqSzFj3t+kPB
Rv0LFnKmrNK4mRNcPdrwwHiaF4dW/yPjNF0sc3dphqVHppE7Ftgl8WeEP6JCgdKsjTqx9YgRegQK
Vh9cnSgaJyq6JaG9UYYKkRfETapa7RbeFkBNAvCGZs+m/RUPh6rmP5YqDNZ+2LASAQOdjg+7kShs
nConMC6K5MECpz6kTKLeORWLXsYBOiLmfxCq9RcxR+HadxX+7tn+A5VxcwWjjXG9+US8FU7Akjrz
5s15+zEOHAXK0lFIS0RWl2wLEf8Tp4QOMhOc+LJoEwNS8SLVcx72nIc5hO4SJR0S6f4fMwdGXOBb
+vb2DGdwUzxtQzr7f4em1Jf9aEcWASh+w5UIWkFDtNcKva8yYtI+f2j4tpeWl00WNiXvDSKunosX
z26J1uZ0QpGWr5rUF4gT/k4FifERPy1ILCesk7aKSDW3UONl1czDkVuwWO/5gbmdd1CzsoQTD2bC
Qtz4og7gdcVxoyCO75Ewkh628QxloptI2iqoFZecBdUgA8qXWuN9XzyuvaSX2bxTe8SZt/+2SYnj
KUKGlUuLRLSVWlgPRqGxr6rp0urpzhxWGrgR17tioOBhVipcINNC2YJ7c8PpKPWUnfH8Oaj/MXaS
IvUVJh5yfuyRrZSVirEXn1JvJX5/iKzl6CnUeT9x/7dFMyiqGGz0NSWrXGZ/QYXvd9t03Ilu3j+y
KdBCktZlSYPWzPgeV3ytLHXUiUjz6XFXvsVCauO6ufwQ4z/s0pfY2eSf0a8dpnXe3x2dwnf2fICd
ysa4PT2MdArFYXXL3MmtTbdji6ncD8vyWwQXuGvzH5vgkyFiUU6q0ZE7xtNQfQ5JtYNowy9MWwH8
xEFML+zdjyAiSnihW04ihVJOCa4fr8SLfH8EZU8pM6pH2pJyXlo78qW9NJHbxEsw3fWbHYyzRQ/y
9SwsO+PQjF0Ae9fIVoYNWLQYRlpoi0+pRJoKJJN4NGiumFaAzTtbRF2BdJPDIrkXe6vZQS+SOp/h
NBwrn8eqhvgdSMI4U3w/YOYluz+w6nFnCR/OsyO4QfX6wJHGbUAyVJ6zG4ZfmBlXnGjdDEXw5MbN
1+YOeA6//bJxR6T0m5qz6pThBWz35StqrpWqOpkSb130qB3ODfMN/Embt9cBbjfSxIiejwej6xtn
xKVxk5fU3eP7Fvrl/LnoQnYYUzOZ92qRs4WcAUuaQfWotR5phIW+zNQ1kf2ZSYSNdcYNnvHTDqNI
EN+zJkrx/0edM0IEyEWX3T5gDz/81xv58gRWNdTXm2DKEddbNUItWNdxuBbVaCbEt/SMMhOCbXmo
opwr3o623ej6klxY4gj7w+JQLIOclz+DC6Tx8mDn3sh7Xvmwsec8ehHfWzj31QRnmggQ2fD9nrHB
I1twQAzh8Ig06UmL/YoSrMKWfOe63PvIy5wPPFe4wevmhbDH6UvGJrfKnHHOQY1oqAOwOH1I/B7l
/T1G/IjpcLpoHAZSTj7YSVoTW43CUYqfPLMMYOHVsgYuzj+dsB+wznO6LVmBe4PejX9oUcjFC6TV
MIDI0fORQSZQzQSrd4gEjM7tg/IFxE6tEAznC4CK1QDLHk3diFNDJukRHG8co/1ZMyznev+Va4gt
7W3PJ3gGwoeQmpCinzC5PT4f60Ljo56xc7LZQhOkVgUbu053v9N5tp+kpRwEKKhllgu8A6Lv62LO
juaD65kPBZL4V8Ohq4iNf896kbvQ/Ek7En5/g5eNKDhzulLivSPFhu7+cv5o6hOObbnLEHUfo155
aePGaC72pGpRzuIuz4BEiL1b6mGuZZtuN90EYKlrYlxkZU2yceyh3h2a5mkyXtaX8VZXPDskn2tQ
a5NfjtiwZQfSLjNVxyZcBWhjWZAbfvH5TpmTK5hgL8ppErwUZNtyeihT09ydRNVssaaTwUSC9tHZ
s2wJb/bJdYHOX4tm0SxiNqbtxmPKVumjqDq3pSnd5oLRUwE45NhFV4q2AZDY6N0OfUTKtktmpbF4
rWeiGt7MKFib1iX5OslkAQy+YGNc3w8SRhYfiGEvoSxNH/NKgvVkDFz6dwsKU5sOVsuVs/kYaWsB
KPhwedOAqog+DCZ8rsuObhbi9p5CY6bktfwHzhqGGHgjiI/2qNZXaHNeBOLUpMOgpmbS3ppDUJlQ
oWwZD/l+1zOecrhvrkALaayvSLAqp6ILP0QUpOY6sw1HUuTP3wdOfUD/HdR8F1gRHMJGpZdbit8W
k/CNmRBXo0Z0D6HcqE3SfjiS318/frcsJOXv5URqyVyINeFWbeyzZv2SCIHIgOXWw3gA5tjFRPV7
OJtUIdPrjUcfV0pyXC/S3Ym1DYP6cciPlG/9cdGd1gNK5TLBKbqTEUqsu5BFN6sHEoBBEW5rk266
fcoKKvU8v0m5UtdfH0zZV3l1TYZh5yO9ebpGwplGui5rYOZv2qpQFzfbx+Mj+oc25TdtKpCnhLdJ
C+V+9yJO1us3VYQp5wr4Oc3X44z9EZF71VjN53qzAL/TOWQWepN6vQAT28cfv2MByWLz+pOmweZo
kbHuJKAR6f2au3o0F1ab1lYmDFCig6d8pDzgmUQKCblafk6y5ry/HBDDId8ysMOxUpnaHJuOY9qo
T1K3o/97hJsybW3Y+riBwSmHd9VHROUScQ3BQcVusT1tzcFzSjO4+u+dkZy5hDSAdUHd1E6i994M
gTQjQq+VR72vex3bn6G9ukjNojMDqqxksvJ3SWJ+LsxyoJIwcwycryJkNgXON4YAg8jn+wh3eH97
sebokI4eSHPV2OnHuwWBsC/dgzn1JjkEULU5veuqVMMatlPqB91I9PXmF+Z16BfxK83HKba5GIQk
SNCmKa7vTNK8NtG2MdOkVqXBIsDJOk/8G8NHFpIS0Eqf7wHXB/nNySRRv3199m+FEB4lXuTK8RoE
4FPbD5Gc1zxLnVEgtym5mXMUWA4Ntb72Ao+XZI4rPu7C9DDxrl5gnvojSmcGr/JFdNLg822SS1F+
8doV5V780AyBhO2o1VQJnytVZdgsP58Nltoa758hBdEoBU4oFnFv3TfSpAm4gQNoe9aKXYY1X9Af
NeajwADntp8WBbfXJHg9JDpMr7JI3lI//I3/yCqIDCCZc8W7mfvlq5AZdwd8eOxGKUIbMVnNTfG+
0NWeZ03hEPFRhlzVJRLs0WbPlNsAmoxiaPjtxTbbVozo25wYq/LKodA1mYU86NJqB3SOiKI62/WH
47rZzsYtuYb0+iaDN5ZrF7tfJ1Z4t5e4waLGyCTAzeSke1fJ3Cn/En8Vjo7aEoTPD7JDjdsUhBZA
j8CpMiMoFBKLSFVcWxdmvZ1Ui4lq6gioRVwGEbjmEMNRIqAT2xh2oIgvfRo+Awu4vwTZkLM5Pu1Y
5z5io2/q7hL6sTib9Avi0B9w4+PgsVpWj38d4D5doAwbrm0U6um+rMYMv7y+0zKWZLtcvK6tiYga
fd2mGDzB++sGB6mfN6/IMoRgjM4dxX8YebWOs2B/eUZfaXDz0qEOJNToks98QCXioCVxNcKjOI7H
eCKkRsnR7leH3cgzrjnByZFIHyhH20SvFQ8om2jMwTxlrZlPg/qU4sDzFYmapLAJmSqBoB+pn96E
Pq4ba/tSF4d4TqoLZmWWM39VwrtIAFK2qHEKqN0AUy8M9Cug+ACDI9NwBSi7tccasXYZOLdwOGuS
LFOZw8p8t83kLVlT4TjrNKgmefTv1Nyq/YnUnDbnAK+BiBVQvT2f+/Xc1TJygzjFf9quvLs7vHJI
399twzB5hUbypCn5j3+a9C8lCjuHhQMozNl6SZB7onNNu6pWPqCK9WKY/3JnSLU8Kqd5P9OrR4Yx
KSdEwCjkJTjOvx2zZfcDrtUdqUjaQkcGs7UrHFpcBW4HMyIZFjVYfnKjhvvwgVIUweOV9c5qbcMy
xaIMlWK21eGE+ZviVJtb22qUYijgj9ac3FuEVdIPVfoLBFbXK5EETmXt33kqapSlV3yoBt/P8n8p
V5vw/HyhKqVAieULVUTYEx36GlwHL9o6Vk7vw998MwtvXEHXZ+3J75v/RNlPMMqaAqjafkNivjRb
cq+5gFQbLWxHHHcUB9gNrvIGkIDnKl9Wt/EofMctUv0nkIHbMZ0lA7SXhfG5oCB9IMfctuYjO368
5gKIWeegpFWXFqYt8uuR6iwNpipD1CQXxeAKmkg295K0h7qb6oYGqGL7WmCaCq87YwW1wGKA1j54
sScJSwUedMBTk0K47pdJ0LH5XAuAAUmc9R+yyHwcv6nzCvfvN4jbkJx/jNAwOw27QhrgWqRDQOCG
N+0a34Y4zN2ZsEy/phkZyEvlEM3bH8XWkos1j5bHNHMdEYU1uPtlubAeallFky6BHQ6VJRQIIMjJ
UQ0XX8FxkKkIrfKfN3z5VMgBGHyiJWRygSFt7p6KTE+jhf4uN8kLUkT3nrn9XoWSFq1AX6nvsTPx
8u+u9SA6cXSTD+1c51R6u32HdqtrPHlfSzyLUkq7ztGAmLSWuRYnZjX8dh40yGfGTNw3cNtBAo2U
4vDO/S2lnyCLALwqseP/7U6upqd5yDOn+rZAkCtPY0I0WtZGPxg9qCtv7qGvMzxSsf9sqEeeZgqo
VLplEfepzwOw7uVXUR1ssvTG+PjPnyEF0lH94x1IxiEKOOVneFysNFGlNaFEZ9j93jmAgtFrFzg3
dBJis5amp/2UUuhPp/5VTWUeUHI3bOKHWi6zhS1HK1xYS9JT01oPVutavkZEjYVw/PLAl5uSEHgD
2areZ5a1C85GgpiEgQqpj+ZFQSphVKP8ZbLcTP/Mx/FHHLYagWDy6VCvPntxGV4C9WHsOCIuvuuM
S1mNJiE/1Ledehneov2kLNk1KEVLxy25tTuFj8Z46BwiawsHrg0H2kSlafF+e9lXpPQauw7Cwf93
h3G8J48rie4SucZGWhKlTNnRW1/LAW++yJKXtd+PFs1vGAhuoPBbOSJSyoDHIrkVmlJWhAQrya+s
Uqj/OC5dDoGai27rX+cpXwv3zkM0AWMPo7hHeSnRWTZXFfncGlXzFst0ZFB9WZZDqBDiVWObw5h8
AuFXP5mv8bEkSAwY4PFmvWuBn6+Cj5PahhQplhVcvNLEofunmdIk/e2lSR4Uc3yp+59eC18LUknB
YHDKzxnywPlZsb/IJhI1Izv98wBzEjxADMUdIGxanOzzmJ5c0dzJL2z9tutlEESTkoHo6JvWWdLN
u+wHqGMx+tLa9OhlPzVQE2PGMgoJTNYo4CBBtB2kTXF2q/I8VPumghLMeiRQRACAZZAUSvILAUOv
CTCKRT9HpgW5JB8/O77ZGuCcOpAwIMz2bHcS3I8Hpzj3945N567wb4J6828fpTawkCsoTjs+5a1C
1IayBH6R5bJKZTe36VHdop96oKBNM5wo/3cs2xq2SFutYJ/PsS/caA/dxvACeMlv//WO7NstBM0B
8WfeZqQIz+nxD0OigM4otqHenWQOzKfhOa5FwVG2hniSP3jTVuPT+IDH75zx8UErJ6E9IYDW/at8
dHEO7xSoq6d/Kyod0ZWHGLXopFGdAjTO9/5W5Uttl3SiOC8dLZ1oaGKVTWJdBcF5nBFEN8VHTO7w
ApkS+4oM9xVS56TAod2kvFjqP2wwIO8pm0giMTbjA+rN2fm59xTpZ5tlzWTALBBPfqwnDsGaIPQA
NVKltLobff+BpUvMFdDD0dFEtq+g5bAVayXWU6Z1dIMpTU98VCwUwqL4eItkxii7JMIcnDsp2pdt
njJYR5mhECUcjmV3aUm/PIjFUdSlKRladHlvKLlOW15li5nQgEAIsX2gna/l9O38kkTuDyt5eqva
Lt0r8ihNc6SnR02b6zJj72hk2UXLQO15Ck1yp65tLKjxrc0Nk1Blq8sZJcP/Sxm4lBdZ45aoNhlr
N3k+37JRhQMv0OLhKVb3AYh2fBqCK/v92CrFfCV4dy5H3LhqA1cPeMtDGq/4eZk9lI4jGwaDHiu6
xtKZ8GRLddZr7479PIzp+IkK8bg5X1+XxdG9ajIiWSWJt9N/7h5xCy3g17O9hlTuJ2y7ar85QIbW
Z3B5GevDywjoxzihzbvFp248Lu98wTeT919dPfIOKe+a1N8z+yiN0GgQl+YD2zuWfoXJVadEAuG2
L4iADeC19U1h4M13lqW8XgGEFTY0pKIsqesJuJw4rD1/KmqBhjkv+OZKlb5wW7dGQCnxL3keATxq
kL1SOPOqOEHx1vv76ltU1Rd+KbgYC1MN7pBC8xd5/87TYjPjGN3Vflh9GDhs0efRcPjhVhwlHfb+
tsF3PlXIuxayiyOujeJTDTonrOzj2PT7NumItXWpfwRz1YNRTVWIqIxhwnBnZptIWnRApKE7xa4i
DmZJlqCG7WlowLIGA4zz91JIgqVwtSugGnS2SJ/XgjuZ6qrvcizljPXbeMUbdNAXYQh8XPaewbE+
irRH1Q+nfpoP6CfSOs6G5kJCRIWSK38QiPV/E4OuMdqIVcBXihE2ofnp9LAr8bSd1Il3EHpD60u7
cXx8fGTDcwsnUYnXdDE+EkvTlKDn3+1j7XjU59yn4G+Sp/M4MrLzAeL4uJjUvvPjXSFN3vvLptc+
/aH0S9XVI7+Za2eKBJy5rRqK0GmvBg25mb/EXIZSH+/CDxBRVg5rjBLGy0TKGE5/4PE0mJUZAb3h
E+2nFXtSmWic3CR8wY1tiPi4vbA1cEE06ZlBJMEdXSsvlLc0VuX1egAZ2hcs+tQ01MNpWOdh9bs4
+3/7Jp7yy464avUdX5zQ4J0JPMXXigZvRhaE3GHAP+zgSt8eXcgr0ZMFHUYHSSZY+jFG/HhL1ten
vtYm+WBTmT5YH6lmUAqprypOiZd6UBulrI2TPYMUdIfOyrqwfsqrugvpH4xzcHVn8JNNXY5FkGoD
4ryBernV2MDm7ZSgMyaaB6olwul+O1bVp4S2x4Jt3GxKR5Ls9du9PKoyHW5bqd2e7cUM7mSvh+mK
tRNMU/Ey+b9wr9NYshn1xiXs+ZyYcM1v6pNLdZIrcP+u5pK3ML6f8piupJLPXfrkT29Z25p1KsqJ
NkR4E+Lq3YlmSA/BDCQb2h978qtSCiuISRIoU6GzSrTqjCWAQJvAVcue9j86FMUpdYuRxsYnuLAY
XpE9JqWfGs3BhMSZPqQDECLNWbDJrYmWTG7NDtkWtkKJLoHQEEwJtmUBfMXQW4SUvT1iLsQo2G6Q
RrXXjYH4R9BnY1T6w2sAHV3w1KmO7C2sl4VwwZYeqdA6tDgrP/jnq2xFKJzQ5ZulT5O3AYj2XkDp
Pbp7WA6y5vp63XBBIrC3YGjMZrrpMBQPfjRCyP2V401PczGOMwBLOZv5vf5D3DariOr9EDCp21hy
YVBgCztdSoMKJK5tCbdvgk1sPTPLdhZWKJhzNwyjuwPNQB43Y/am8eSkSDJBnJ78asB+SZqRJKV2
apoOYRFZO0blK+ymFdMA8f0aCPZutdFOr8Z9fqvqAeKZ5XtFGhFAeX91P0meX16k2m5QKZ872mmy
bVISWgcsAWUIUpzZu0LKpCZ+o9EqsfM23Dhh1mPRuwaMp/ynuqFfKxYnU+1AI5eDrIeUD5YtgvTY
0uZetBM1S6TzyFESFDgTfHRfgpupn9VRyRnZrJNEcvfycWeynMzQ4r846idNPwwPpta1HKzY78oi
M17gTqrDUXywJ0jXqS6FmQ4fGvpPgRRss4HpsQZ1J+WGcLgbol49yMBpHkt6sQrDHWqtF+U1F3lo
o+W9ukBCx+Y5L83vlLE1i0v5GzKbpr1KbhL+sFIgcceW0uT4tQnLWOq6Hsc3piFEuo6AeiJFXr5U
3C9isbmjc5xyGvIj3mhf0lhAQUFbdzENP+MH1CFPoxzjhfrwJrEIk9z2Qp7PPcbmloQmDfQ31fJj
G0vK3Hclben45HLqvYnAzzc9KfUxt5m7h1EOWNEx6gDn2A0wECksnxJQVjRoSC3a1+yk59kpTr8F
1vIZcVrUVIEEqCpwfqsqNhBRySwW/3KGd6DR+LWbVsF/Ct9j0A7ljsn4KDj1a89GLr1ZLWveJYCd
iqWIDivVF3qNJVTmL9mf+6t8CAzu8ET/aBM9y9bgCW3M+hm9D6tbK0zZiy+ZaTh3qrEtnI2bJbGV
70ovzVUnNYluDnHIvLtu7O0hO959GAz0R0Rlw/uzssKCjruTXAPyyMBP7fb/BaFzGRngiYQtMo+g
8HWqGFw4j2BUBsKikjLYTHFcvwLl7lkuXDIJ9QD2oUHMKLrpr6lvANG50ZMUg3jgsGiZl8OKrbiY
hjt30Fjsw8+VqWbxnr9YGL6N5hc1TPsyghZDMKsQ2gCuv+tF8aeBTtXqrS3tc1CmExUc/X+5DFTV
UQnSGSAgE4KYo4X7UpwHQR/GBdrdkcTOScgpOjX4ATUZwzuxjDtobZVa5KepbBNln0PdJ8GJzsTK
MfBrvSgMhBy8zdwv1wQBYkxNxTCfco8XeLQeg6EzpMd7MIbSROLrEkWt8RImkSR0SbhhaIuwiNQS
CGSpiQVUDmkHU/0Wh1Hwb/xHT2AGZc9lk1eNtdOv0PHOruOzcRHNhCQe45t459xjORQWd/XCkR6S
Y2OPAKKryWr1pKBF6OfSjBYQUEZeRaGoIEGZBt/TrCMkZA3NdcWgMdIDqLKT9z+S0WFCF+c0Wyvn
Y9OS4W1DPYypNQTM2uxP8IxFTlohX7k6B5DciC2ro0Wg1ZkUbyBv5HKtQ73kw8p+QhskDh/dpHLu
fjtiDRqcQjf6LBXskfqQc3oH5AYWiL+ZCtStFnoIAhJMnWeb32atY9lCwTgPu4J0xopZJt8jausd
jcPEOgR+8QxPuueQpeKw2pw3Qajyh2YhRSSEeA/b0yTH3mffCekXNhk8SxNnAdF/+RhJ6AxCBVIY
+qGcQQDJGTPfPWkkY3Da0x7VOpvlbgcZ5KuDwUee8nBpX7jbMOtxnMYgCrBn/BsJ+nASpLPF4k7N
FaUN358lmz0KU+uYzKE9bFOKOeQNqXLW37VA6Cm91lfbSdFHaRMFFFlXWo1r37Y53OAkArIpnwzj
GlfmqHet883MZbrRhusgIYSSIe8vPHm2TBhSncpe+sd4b8jJUf5s4bSBPcWIdb8nRWDQidHTX74K
e8BeFfcqHgYW/9On1gidAp3tVrkfamAo/mf5RywxVpcoh1rdEbt9AxuVrvdTaRwYdndZ9x2Orfjp
Sz/bhSiRw6p8yxVd0r+VA4rsAUldXrPtA0fbmYrMPABYWPCNr0eNwDTL4IrVb/tvFDQnBvXXb4EZ
HIrBzWpTr38q2zZHDUbKjTvbMQNrGgaAo6i/gKnwqPJdJWK/aZ2Kird5LXFQvc3E/S8mwYfZjYMX
3SFTrSfCkHZomdOvxcVtcaouQxrrfzFQYc/fasuyKcChrp/oo/GfKeGpB2Qt2xQtG74TU+oy5IWy
KpVC6mJOgJ0wHFx/8FD4MJmGZgE5hJsztTkEZemKdDsUW627ouwECl4WoG5fSlwKQh8PNJlUQfIe
ftd3AO/csvc5sJ2QOymopywqV5hYm2HtDCF9SZF3MuUlcB6osyBrmEqIFr7UMn0OS67LAVXBgOlR
GbXuTtmQ3BWhAQOzLs00dFP6focqoj8VuOBP++/4NlYAhNj40w78kscdY2fC8tKX8A96CyX86qtq
12ka0fzY7PfIkjWxQbfBhi78/6XBYftV0ZqP2T/r4DXurlLklo32GXoexUv+tdN7zK8FL0AUJq70
kz7yv2Kl7cUEJsxNnHjC64xgMZnLEhbD7l6NnKax4+OjjE0egFyEcosw9OeOzDSTt0yEd6fBdkHK
CO1kcoDr2aezEIVEafp9T91ckjcp+l1owQUYsMZqBsyzKqZoFJ3VpCuZk2eclgNcpL5N0ihJ26GZ
s4SSEkoJdDlKSrXBNMtTR9zZY91rz9HTxqIxmNduStMaNjqOrvbtFv0WnnAf8pKVpgtyxWZbN4Gq
ZteuuEQkiHJ7bV1iPHqLVuori1FSvTXyo1Vtssh0Ed7c7XzijL0+o5y3GwfIkVXp142y2w6JfjEJ
fLGzFS61P/7iX5ndalBNG1VHteMIlxwD7kes8RX4KlVsZPfEdfiWP67esmrzsS/b0XmyjfZLiu2F
0/P5M6VMibWx9JXX0RVlTcFLCvw1A2SSMvo4Q1Y46RzlNGntoPgTr2f/QH6mCBtm3+btA9jGkNng
SGlmmVexUwOexeRe/c3lV0DBNUj2dA+Mfmuxf78A9AIIY084HNx4w2/l6CJxr04RCaCmb0jzTp/s
4GLcxnTl1VMRYcEvBt1H76sSUv7HFTttoIOMag2BSFLjdW0LJdU3Dmwt+BwPgihZHvDJC22XHJY4
1lLh1hLTIRIQTJw5AZ7VzTzEDvQzOMx6iQd8rp26UzD2UN/4ghorfBTnkYP/Nvm0orwPDxVpTn3M
AUZq6DuNfQv0ktrMkgmU+Az+WzXn1lj0XGHRGTAHjbhoI9eByIfibl4NVnqh8A0GIiCuYfIGETQ1
AeQlkmbiiiUowy/LdBiRGIXNJhnVB9z1APw+sEYZOWMiYEbGae3sXnPqsg3wBrdHqMAmZF1Kle+d
ziGYgZDbBNMh/p2FD0qIl1Ebl9hKNxrH83CNBQ0TO6Oil0vYU86yLADchIQUe8105gBd/enkbJfE
kPHP1ywPhzRcCFw+fhBn/pKjZqM8X7RpNEHVsSPFFPS4Gk9lhin8S9uhNAFTeTBIB0du3Bh1VjJo
5ZrGekuLD1g1gYXeKx6NZIvTr9/m0EQst05+Zy64kY7WfxI7KVWY8j/Q9K6QqOKPPuHevKFmxb3N
enA89WPs61GLcmATBEQmppvjhN2WqvW0i2Z82uNWvrc8Q7jv8d0q5I2K+AkLNd9JB9UX+Nhi5JoY
J1hnaa8bJ9i2ByngZZoiLAeslBTlZcfbmJNlLTZuI8aHRTzMKfCSTQpvXBKZMq8ACgO2xo4I5Ov7
QyPup0yYrEy6UgnmRQpZ6YgWSP3loYy/IYaH61bVytMINPekuIV6F1h5JcwKX43Z9ZvWovsIQbpN
SFwpaTmmLmqWECHbhnbWrq41pF8oTlp4PFgplNMs9unYOZ7rT8yyAdI1q6fFqWLl3xRIZl+vgzFr
ELf9SDkXMOg9ID6kWxvUvwxg8UJHlNKCvQOg/UpF87hLeHkbthVJMxmt6NuclHI4m0vZ5+Ybg8lS
xSGboVc0L12rDqFu0yxqUbJsWQkydLQhl8pYQeEnOMD37ZdDgURP6JP9wXKktjIX+OfPLxjLHC+t
TAFfN9XGnYFj8RvjarY6lW3w5h7Qt6ZdzWDmgln42d1a2BGnDETtswnkHe+3p5SVbQ41ME1A9arq
ZKVE3GMtG05PAxIgkMx4pmMuylbgJhSzxMyqvdZHKToWEBLoFS5K3CjpbCY9XpRAAeya0LngmcI4
U46miE29E+BCP4K3pl0Ot0ahsTNdf+Z2FuHbdu9MKvCnXFm863VO8bEHrjQB4AX7yuUJIkq+NNqP
T8bfO3djTtBBEkTcN7vHfeRDqtUBcsQY4l+DtKabKt/F0b3brOv6oDAkObCu/mf6TXHqMrETgnXy
0T6LTlKoSBXvIeLabcpPrfvgoZoZl2ddwyKm939Zc9Q9hS4O6MepNcY5+25fWjB1zSyedmzhV8ka
lD+6rn5zPRb3NclJopbuAP1yD6A88cITbqAqIiQ4nY/e9X6h+J3oOqXzFM7kVKR6KAbpuk1d72a1
dz/wOrSnrX9PV56s8Rb2h3kC5u7MXtEVAosCUKe13uQdVXWDhvydWEfGWAu3wVBCV/ZJMAb5zTuY
n0aYw7BLy4Rgc1f2YqtiFt0vObJrbNJJ1Y+vPbaxJzsRbOMz0fbqOU6svL0gUrkwdE0gkXOT4ibk
pak4S9pW0LS+1RWX1gAp9uXdhgcTY1rrFoyjNkAAYG9fus9qBoQ+metxl6OyqNKif6xLF2Gv2oVA
e0857I9VnqtIpTiM04+3rQhgK63SsE+9MqlUt2KEA++aawY976uMdHNH/aBo3BoSEl4L5ZvaFAL0
/dH1BrPmIsZ045N6xA76gpjQ5L2c2xETcQKzn9rFkcoHs1y3dX/HQu/5bbNduZlAt8vj/xpJjX2d
KIDBl8VccHCa/XU/9QCmZRnsrtNvzTSxy9qk0LIf8g1ki2Y3GYNpxCtQZZ1EZGgcQ8CC5RJ8aYD5
+KqrryqH8sGkbAqVm1weQsCDhXbqXERq2ezaiERBl5mCzqbiJb6zgusayf1AVlQceD2UDG4b4bEW
dOPTWw8hQX05kkZMxNPmyRhiiqW4GwrtmfSfNtHR0X+Z60tJrJHHslqjZ2TmghG04DSZZzmZJBC1
WdnqE6L1r0XrJ+5oZGsI+GrpBYI9DYBQKOI+UT9QDLkV/iicktCF9z+sf1svGgSHR2RgLMnNaCWz
M+ocWQ6dKk6ANJchK/4ZeDm2hXbWcq+9cyiHslVHfRCwbh6zhA59UBXowCdrd4f9+fnc0vp8La42
S5QQ/MleaZvg1k6DrSs9cKF+euBP0QkYj3xpFXqKex1k0PlQW8HAcq2U8ZEYFzCmxhf2CjAJTnNA
V8nhWn8ColQHbkpE/UNjyNzeIET7Qf2gnDM1hwlVUGUK8NfW+VGK68VDnpWwUlZGT4LzA+jQ2LRr
QaUYtW2P8zL8ywZCiz8CnxAshOJRp7tE0yMVTg3NR0QZhz57sWXax6Rxn6W7NMDQMw4zodMCqXmd
JOYugWPvh9Kx2NroUJz0QC9s1q2heLDmgdjs84PKCHwCQTYhAp5X56Iwdal+6m7Cn/5t08Wf6aW2
54k9qcIXasSpuampral6d0/Qht+4fE47NOO36FGzpluOOJFJqw+E0f2fr4eghdDtEjre5m/hDpey
0d5adStS/2P/MRu/h8Av0h8WKu07W2abqqtmxZpPABtflZh219O0J+KfQmOYBiaDo27AXA5YSsLm
Gh4N3ine80I8d03IRdT5u8Y7ui9CYPY40+XuldaNlfTrlpOmyYZlBu02B5mu8hBVNb258No1YKJa
2fN9xzAOTKhuen3fDPsSGwVny/W0StD9JBW6prgmUkZVMHQ5/oZiIxVe+SsyVVCPkHllqpPF2AAg
vILErnBQw7l/dXAY6WyL6iEoWq3utCCiG79ZTerLjohg1zaMXAGzeWcCWvM0KPmhdcQWfhTvvCYR
ut4HIAr+yoWXPKfy0fnT34JOYaSde2wd3USkJgKNAc1mz2uqpDh2Qmqp6IUMpbITjaa3hNi5kAHA
+R5tY66TcKCeYfgD82nUNCrrax06b8K/i2akiVD9PNzv6D2A5dEbpYf6NQaEkGVmg3x6YviW85GN
rz7pDeZN4Nk+cMuaMRvEzO4Gzys2qdm31AfBuYnGME8JAkyYHGrf4QCabFGTqpK6fdcbrHPXtWQt
BzV5rsYuxHiS5i5jTUkYq3MGzBjzhgqVA0nX1VU8k4uorGDE/bPGb4YDivugXuoTTUs6cVqTwvpm
uGBxINwPZJfE5f4Cxkpvzd+FjEUf+jPA5neeTGoumqrNdTC2GqVTy2Uq+3SmU2m0IvkktbW4Cyin
fvF1aplh+pZnecP/AhWhBs0G5OstqCR+5IXgh9HyeJdybEG3rhpzRfAB7uIRU2ZxwUOVHtI/x0UY
9CGZKmRM1/cUxVD9CC2m6Nf66XYg2pRetX5HzifqxraxGVt1vEIX0av89PVKlNSVnDsW1PAW1cBZ
qdVd8uaWLksIHtPFL7z/cF5LdM6SUGAA23yfbgG4gCOEfgFxme+oQVQTIu94IxnxAJZ1Qnkjy13+
pRQvuQhE95qtTN2acCsn7EzPER2DMp31k6h34m/WVHuQs/nAYoEYIMWMFMxjq9swrrmCnYQqRa3x
dkLlyDsfIRgVFla8lx3KKy1SDKDYO1QeWskbvC+XPjspQme1Wa82gnXIvIuVAY0Pzh7ATECklzdi
E/debwmXdOPHvsNAjIahBHvl935yzDQxypS84R8jbfNG7ZFFHHdkDR5fbvk6W5IUQFNEdWI0u6ig
1qd1FkXs2TPzqQLc0gTdjuVkEkLTCj0xI5YTTESLv0agcCsodn9g3v1dfJ9YD7j5QDyb3LowdtZI
8Y+nUjqBv0nc7u1Trtw0lHi1jmvrEj6jUGeI1bsOyzyVUoa9yZgQYmhxit1fksSmc2MeEQX3iEIm
zOm/9qNNaSDqBBSw9q1Wzw7B9A21U1stWZZCEyUXY/jYjy7yZVUaLJmYars97eKo9a5LpSkKmJjG
2rTSfg707O5zLPJkqrPllRfNvexIMUrTFbGsyLpBkttHXI5BXNinyw42jLh7NXPkqasaX6extc1s
AZBoJ6rtCUymbgKBQMg73mifbYkjk8KJVtODSA5LtukC8EWTNlbsrG3r12TyAMC6yZlDUJAL6dck
lLSi85HKsKH/gG61W+df7dTD0Xom/vhYHBVKG33NhKnqf9bLP4fzMNg6bMKYlk4jpd6d5KJ4rXuZ
Pr58lClhSg+LWWKCmh4cGqGdEheVNsv7/nmjDHB+Ls+B1Mn2qeIMKGzQL+HcEUgZNIs2nhM11tSW
DkXEGiaohkrM4xk2fxIB1zEXq5cSzfcdTT1ZR/G+gQHVH4T2We9RM9k5RpO7GbhiTOsq26WQe64q
1/zurHnGkhaTmVs3j0xpVq1iPc4KwMvO4pbcCT5/wTphaHT/W3iW+fgvMCuXVUlqZbdT5135UAFc
2jKY8Dl4cUnGfx0R8CunU/heP+Y1vNHJrpJZ65ABThpyFAFaWgEfNlL/asDPFa7bs1UaKYjr6j/J
HT8NjQokrm2LG3CimBZHBy9piLlDjiwsr0PrJiX1kxVD3XHo6SiqgDpzYHMXxSeNAPzYg345UhLI
FmergethzrO4Y/ERwXkEw7YwzKhP0VAU0u+LB97/pI0QIl88RZnq176SI7/7KBf+jEj8rzB4LurE
yu8E6NQ1iVd4VkCVFpcjT0Qt6zseKmaDFahMyPEFoMclAV66Qxqiz9IiKBB0pT6gK0g9vzBvMkwA
17rI8UZOLJpqK4+YkCmoIelWTdZLCP39Md4abxptEAt+iWpHplvi6ZJDa9S26g9QhIQCwyDUFzOj
BxUl9Kyk5LmLXMcu4326Y3R1OGun6Sl3HvWuLgF3cwusKT5ysJZCe0+J4KgJsBbGG4NtLW+XfVdT
FmG3gZBHNJO6HEfBpa95zXmCy0E7k4gllWobfj1vMRH69ucs4XhzLF5raowm1a0jGacg75Dk07+t
WsVaybnAAW7wU+gDDR9LumDVRmQ47YRZ4sbgPtzSubGN4BYyfChs/ukf36yHtv3VzW2sey99g2GK
9c+rW/NmhEPxM/mdxjfRiyODbBlISaPHsr62l8+TF7ZlteEGur1dvjKEIvUcusBJZSazv2usf9+3
1R35y0FvcT2zlv8CYwuwSdLCBoAujYLjkzxlh+vKth3FfhvHuX9FwiUHQvRA5yn6GNzU43mSk92d
76vshCJh709TxARPutoUH+YqGCG0fNLUVLhKuAi8EGdjDVFQSMSCjwxa9KGmqIBpYmM1I5WyimKV
H2o32BBnhzRnJo0VPWhGG4rtdpOc/RQwxPygL63Kb92eP1u8H7C2etbUtz5Zi+KUrHLqe0e2WSJr
02sStZ5du1m1hLU+EURl1++AqQYgWzetCJbxfUb5xXZeRG8iW7UUIatBLsbUZ8YzYDbprjSPS70F
qDVNKjgCBJROKC4KP1kRI/D3SklFiQFZziMAF6j4N4YJjVdY+ZYm5L25r3fhQwXsb8N9Jlrpa+d2
nrCTUUbmaXp7yhYKNq2dTUtj7lthcaN96Khl1OzLS4ucT7kRHqYREY7qdXRpJOeCEytWFvLqURVg
nv/hkZJh9tcr+7DvK53xqMGDmQpsoXw6UutxNEt30GsTDSRvAUo9akjiFgo9QLNmnU+pECW9B1o0
ufMMLAJIsYE25tyl3iRiWx1UAxkNU+gs/79JNtur/Dgg99YFyPNmYY0a5hH/m/9zlGjX/lXZ9P4s
CmrihyQF+SzvHng2O8TP0ctD4tbQhyeyOvk63WCTcpeljvNxlmpDM11tkcppT7OLzk2/FZ0xU79K
WIMJhLgFXEJokhohWO5viFaqr1bf1asU5kA9ZAvuLE+UnBpEuRbDXRfZ5AuHq3zE7XRQ4/7RvXFL
eYHy6reQsBcQsFI+NteiXlMGpOTUPptt9BonsHu38sdLB4Vg+ztDWzk9zrliQl5ErfZ7Jxe4iFXD
WVR0LnhMqqLPjxgyh+lEmU5oSxcg+sbMng4E+CIKPusQ9ahPlCXVKKPnIHo3E+kj5wsLIYAqYIhB
zpxbzj8//Bj+EeO/S00Ymj8ftnDdykqkyCURGHU8lnYw9QbuDMscdFxTlZPbM6gofZ7avNt8V0/h
wKxhj8eCke29wB9XE6OdxZlLQ4IoEJ3ngB4q4iYxcp5URnIN0SofQDJu5z9q+S22v/CiFH1+055W
SXkMSqM7jnbS6gZCybUJoryrIVh51g4eWAFyhAocaiGnj671+ypHi+PmVysBkypfi0xbhDbl68Pa
v+AqRX3IxR3JE212KPK3wkrw6dtzlMSz2lQ2od0LkT73oMLJYH8Gv+hebJ8mgBn68RIEhMLe7fvP
4o41hJ5qGD2ArO48pJZ3RgMeUkoXS7Sa5Ii0Wlnqjt2pYFojw5OQ+2StfO8IwVMV6mhqKQlTUVrq
4udgPcVfpTB05ZF82X+chQQw2Oh2a1P6t2pnlzfRSVPLKqMRE6hfKSbAqHy1V1+fJQjaZNZUgm5L
dwDMRlkjj7ILnO3gTcTgxHzr3h5X7XU5HTMiX8FOsVPcWvvybJSo9cxlUR/Ob2Ft/L9R79rZq5ns
tCcnmlp0eVQ6HntGU8ygd4E537gyIrTOdDvLf9npy8aU9F3GdYpP+LqIeZIg0i7Sx6fMHckMs7yA
oLsL+kZ0ivdajHRBawXeki2ERTgf3yF90lJf9MTgnjDI/rMNRbAaUHBeU0vEa0swMeYPq/H0Um6U
fGPsxvXD8f3/r0S3GgrafVDsv7T458AIsRtmW6G1JLQjewk9rjaaGTZ4o1t7W2Im76PO9bnQPeTu
Zt1szc1Q4N8HXK3l5lojtL0NY4uf+MrOhqtmMByilw6dGT8W+e6ZKXxPHdyc3pPtDwjlM41jyKCm
vfWD3PIbfaZg+szKEloZpMqT4jE4YkXP/uatC2qGOIzqYXwWeacCufqK4qCaXr/PAj80hHh9/UtQ
iyPW4Ys1Cw9WjNhWAOd4vfV6jbtdYYFzFAD5RzEkOXzstx7r+XTIs4O7lIb1Q983890bklGZdcHD
h4kGrvByzC70Tx5bKM4k2nwbXJbIHdHiJ84m+jw3vAQduFJuHv1zFrql38HBA+B4nVnwUe+i2zg3
QbEg61JOYvUqLXH+6LpWyV6Z1bXszqUWdSRK0h0VKAgvJFnxlbd7MLWmCGm1EEOOG9El1phrRwaO
lSg2c2DLrx7DsXg4c3qyAn28aIGb4cL0jL+681daSrX2gdQF/I9F8PRc1b16WnYTpdOoYu9SH78+
FIrZGBHm40eKrmGECKuInCA4fAK4N+lkCucO7Abgoc3Od/nJ+ZrmvbGEpmTKcUwjisXwc1c2KQZw
hOLSSrnGJWaCLD6C1A30Xmi37fJQ/AyWGBYeVq4UqjpWzAhle8lEmY6xZgr8zMFRWMvOTROif8DW
8+7R2TXUuH9bSCSdV0gk8zhyBjIfcwXZg2svHoOgmz/WCPfK57y2zxDMQx56xqdnQDrGr7DC507C
QF2RMyQESI33umTo1tfVMDDDffth7ZURro+PoufpDFPoO4UOuvbRjAZbeQZyD8ube2XyfMNd6GaA
kcnN0UxrJuFZzxTnHidJ25V6cVAqPHyEe1Vg26omNOkHLI6sCq56yXXhJiacjq7/goieCdgdjTS/
s61RWt6qhwi04vh5l0VS5cmaXDQ7T5+XenP3Cma3OBIrDPEs69jRL3sWGXNvO+EOkykUfguH22gW
9EJHTY9MJFCuuuvm7TF5G4ONKyF9BsRrNxj6s2Uh4dmCmFteGXGuumyJBRw6iQHQNnHUaWfiGEfs
YFBGjrwaD9mP3eE9GSuOutWaEOFHRMAwNGhM2LXa25wp7cOQnwUpTqFEvV8Splowib9hHC766Q0G
ssQNDP0NHiu9X1ajJQgDvUyzr6xaOopdGglGbtxOsL19LnQianMr7wKaXnrX6uJJIJ9wc6csP8M+
aFDhV1zmlLh5fLZylsXfRvFxeJ5mLF260QOLf7a7KYxiT30Eq0RvvEmcI2exvgX0qRl8ep1XYpi6
hUQipPfS4LZnGeArYF7Fz+Zw9uLC0QXoh+enaeC2yRCr4zSNWo6Y0ZG5ZVnpeF6EtpC1bjIEwiQH
7UUOK3R3b9Ps2QgWYzyc7ZP/jV7gFBqL/51HxhobqMycoHDvB/+j1B28BZnaqfa6i0FHUi+V4Kg8
lpuEYDzuawcvFMOEHiMqM9qUxJpYK5OBWDnytRYL+2eXAoD8Jhg9c2iyzfVsPpWWk1n3ruWKmMjd
zJAEfNAMjm/1RF8oohUrUcU4qyPQUbuQQNzfCYzZP1ST6TA/xzoXna3fFy8T+EpbPodRds+wc50j
ammfYPiEEwe9nnoBBroAvJdslMRCms7T+M1G2gDNPd4svxOu3tHY0Qvu0jI4Paxt3ZqUtRWmv8j0
iDCodMR2P1PctQ4lWfcubUboE+DQgcGHL5Sc2xhwb5miSBOekV/kFho3+lPjYMGL3yMx/VbrH3KY
cWcmuvI1WuHltCNSvZcPCqoCEVrFeqA0QBv+hb0bGUZxje0pUC9fx4Sd8datTonD8pvfRmBLT/Ur
1gM5qWTp5Uc3V1uYL5SpEN0N9MF9P8rm1pRdIrhDprPXW/45DWHqGubxrU9BqHFiieW95hl3ztzI
B4sNfNfxVexbPdqtvHzrpcPIhOA5V9WAUmOy7hlSv1Vj1bcz9cI8NPd38eCInDNwL2rE+vKN/jdM
n/seTH6ZlYV2fi1moi+KrNi+ZtbQGEmYJ9OlGXy+17OTUC7BJOUCX8YESvsG2JxPr69WJ3bbwbMt
cmApJZy/mj1/JpWiTokLQ4WBV+rza6O9MgsBx2d7jMhBummya5o4kZHHJEIV04S2WJsX6mN+clFd
+jPDsATNNzHRGxfCZES9U8p/5jBKRs7gcX2lX5a3yqbu6cs9sKlwxXewjPnYxCO86rcaiF/J0omr
y4dTzxdG+u6/gzgxbqbYGZ8dqdcN0iDNmqzGBHGr24bki02oeXDLFoNxLdhPVeuaeyULRfV8/Ozq
dmGf8hjO6TyXC1B0A9dFzagf5K6/lWoww5oMrfUn1+cOIJmk/KVpFwCJZcvAwujpnj6w7lh49xgN
OQ0V04K2EUW6Zv0onyiEzlh7Fj+p983Aj1TUBfALjZHVv7qi3ZmQ+gBwbvR1PItih9p57GXbnhhp
0CGPu8XS2IkhK2zKb5fdqh/IQQ7nCIY7mNug2s8Ig04vs3ECv9T1aVWG7z7n4vqyJ7ixTwCzZR2z
/joDdN/t8681ZEUF0BhQrlHes4+MukSRJ8NybckY0ec93Wt6L1PJb6yDbVRl44lOGkl5u4p19+YQ
f0jzbtSs0hZNHT2ETuITZABCHqNu0/1CAaTO3CrXkETkwJkgSEpKdm1nJlwB+W1XdUOvSj1W+P1N
scEhKq6BCFf2uh/nHHnp8vVwr+JH3XoRlSxR8nAzfc0LTJQNdzNWQt+m8YossrcXdr8DmUwFsksJ
SQeELJ+NBNZ/kagTYs0ta1UpbU6QHMWPpAe//YkvZo81OMahJwGhJp6I7c3LUMV6IEO9ycbinD+g
cHZz4gSPSBTfla3YpcFdjEm7Kn7NFZfoLHQoDlfz0FUFiPGvWiMGSuddgy+x/EKenTBCErbs7viS
2ffCkXeZ4aONa51CYktSFpgjDtoJUarWBKuoeD2TYZ7UbyPtIK+aFWrrMcmREffb4lRrz4QJmu6R
mxvKa805ijrskRH8pFzfvFJmUWvwavua613XdbDi4khG1ZSCUv8RXgouyw7c7E1ovJtVk9xUHMex
AkuGeeWNwdGTu5XnI/EjVBcLTHZ1BGKLW0SfOTird6h2sMsA7PdDnYe06I5yrU0FttDL9+Vd9xp1
0EE91R7sQMtwRQ+5KJ5v7MyB3tlihf6C55W2JzqrbaBkFS5Wqjak5HT7AJsB+jQD+GeZe9+dK1a/
OWzak8jUst1keKh6fEVQrbfaqu3I550CPAdZxzWBEfxv7ZstLq+cGspiLweQKZUOzNgV2HQM2QGc
L65H9uGoGiwLmcH8uA7VJQ/vAjYQzxQb2Uf7OAxuuQOLwfkhwdYGaDczFPeBYp+c+cYD6ukaQ+Y2
PvTOu1tUJUfKvygzxf+VBKQOxqXDRz9bCv4MHdjsLt3gu+BsWzeP1PmBfh7sagdCpIrEuS3+0q4L
AoEbCqCU/y6Qt5sXz7CoeWfzC7EMHxEI2lRtZSTQaveAS19AzG48ADauMtk39O42k3b3fdzAfH5h
jygpMZodjt7C7gYY3j/GN3RgZMH9ORo42Dq51len3y7GQFhgLRsdfmrwPHTPv7mvFctQ8TdT6VkN
DdaGnVvQvQigLpuhdK7kmzIJjPHrZwdqipjVw0zDgEMVv9QNaFVojvtuX9T5dA2XAuwB8JMshT9W
DlLctDU8Zfanm31kyDbVP0e7UoAkjk5QKsvsEfQD/gwRZlFPItfvMTbptyIbOWCFvJsxvaDHJtTI
m0hJkexr2Te+QD0n4xg2HZw5p1EJPZ4a/xJBmWT0iGOqRqA7gWc46M8BPk0QuwbL9wgr9JKZt2sV
q24+wl2WhExR0kH10RMLVesEHmm8lzB/YTwMa/B0x2Myw2Cn0qdsClenzIb+WZcJLwYv6fvn388j
4w7gpSN0W/fQdmpXs8qlaA0tgBZfwpJ+O8Jfa824yVyLxb/Q3Jl9kwu8PSeRF2VKstcvZpqMTV2+
G5gNuja0hyEkWi93drfoJt8TSmSAQXCEPYuFBbyfMF73FYEx/uftA7ABkX3wy+lS1EEhgKgL5H1v
CLn1T3q6+gGVDbGt49KXItISbm27QOZO1AmpMdE3Fpc8978OhguFtpAGjLFUjSiqjCrW4btVEVAw
VibQc2pgdW04vkPQAwhqxDwyaJh+x4BzR/h3YxwQ7aEnGnh7RVIIgLdMDdtwROfkJt+f7/1BhqUR
eCTHagQqguMCSox8aqIPeMFRS7Nlo6ooW6JfQsug4PBuQkaYfpokzIRZNkMb9L4emmg9GDEDvf0R
ChRm67ECClNCqj/tkXKPoDLlroPPyPS/3eD+OzZKI4sncaSVd9K0pGyHygPp7wSLhqwoXNM/LqN0
3iE/Jfy0PIAhLMXKzzg9VtDXKx3QT4b08aj7QyQXfbboLd8mgoWMKS2fIzVBzGb09uQqzDWNVkkl
IhzozCJaaDt0Se+5e6GWHkuMuRYKTfQU2+vE9VWDqhOJVBp1T7f9tLOJZC/15csw7dcLEveNccoz
cygPa2LeUEKZJdin9KvA1HHqNv/QXPnzc8b+TnJUQa09SZzCew4AuQS62R6uk8ukFSvvFSmFGQR5
Z+HcsFcCZ6f8/f/mMC7ciSwNQ37t0wkvhZGpAUBoaEVc8u/pNKg7s3Cjd4c3jIbjYMHdchulkDEU
yuZOWeD6N+791McWnC0QowPGSCYdt/i6kJVUR8sxY0F5p2OIzzJ9y0HW0cYNhfOY1fEcOCXN8aEf
SFe9/aEyeg4HFhvNsULgI3XzE2txceWwXuVb75nqNXinlJI1V1JOu8OgAE9oEgGfdjEO3IW8ZCMB
4wVPljVCz+lAl4RpKjrE4iaZypSlmraonHPmX29DGCQ8fjp+qE/vJe3mp5OcGVzB1VOhfj4gej6+
xdBoy0eFtq1T9BYfRcW3iz64WBqbSUVBROXMXJPacgLKjZ029xJqFp7YY/A2PSMH3l+lmseOD/R0
bB1KqzMY5ODF6y7G4PKNgexGCI8QZ4d+jr+M/vfER+q8d7jHgYD6xFRLvAW8b0/TMp8bWLWF059s
XbWVAU2SGdqyfiG+lFGEjMYvrbnmqAMbw4whgxbwMZWSUoWV0kaD7Y7xixQnQ4Ve6jWSltCx3xvQ
Orz2mqm95Wr6pgPhJWQBuUFA0l0azOFdaiCu8gR13uHRVQ8+bVGzustSH4xemt2lXlkqiL2HN/od
Zc/LxZHAU2dwX5ruNlhHceW+T7D5R6DmCuz5uuo4ckw5oGD57jOEoWrXU0GZ6/GrZrgyn+5qyKPQ
/PZ7ZG7tLszykVJxN395zm54Kiffh+SsjJX7hWapvIsv8dErk75IXsfUmsT/3kz7cV6+qSbOJohC
k30J2dZE/R6OSEPrZtiqsYb8JePi+c9YXErGD7AVR5dbSvF2crTZxSEPntlWErUKgJPQKarn/dMt
yleraXIjTzzyMR1pIwObJU4RO+wHb1k3hz6/fP9KSZoz9rZymkq+54WjNwczvYN1Cq6WQH0VGU9T
5ncwd4B8o16dng6G5a2CkRHJxi/a6WlM5SkOVomOW6VgHShtIvzCbpzQONP7ZBV6Rsv9V8+3PuZd
cwfDnIY3GSMhCOfl+IuTBueoEmo+s1lq6I/IVdPLf9jo6Idt8sKNwdMvAcrMvsHAAkYPu7YBETHH
CrrrTMvYT5qO8YuvpPvvQJVwRy9+RjX10X8jpAR8MBXWncj7Lgj0AZMxLr8Vahm4MG1yi1GCejZr
5fiRbXdw/VnzSlSI6K6EAW7s8OpExylMlLkXEfwsSh7Y2TJDQ2NVshx8H5Fv+A7aCOxwHmgbjXFk
K2HLsxMSXC3YzbxEHkZ8+966VPVQespGpahs/9lV0bJ4BxFRN4jy79Jh7mYuowi2bn3Q/nMdgSMO
K75NrnUnc+oDESWXdLsNMwUz4ySUKB7cqLSNWJ52M83DpsskUyaBen+1UqXgoc5rBH7uN8Q9VoJW
mvD/Oyg8mZws8aBzIoHBSE28FLJylW1qq0aaM/n3Wx0mC2RGKuU2pW1xuz1AtyYtsZXtCKJYsYNz
8KnDjikfPWHZkHFeUXGD9z1xGGCXokn3IQq3oA++QB7tTuJv23Rq/h8wxTDYHCYaNsKMJCJdEM+/
xFBk1Ekn7cChoZwa+pCQBOcdyWjauv1COXsuTTwjkA0aRZgr6Vd8PqCoumjhqVOuKAN3snT7cvX5
sel/sxe2VYqqBUoD/d6xrS3Q76DC7Dv5MXmyAi0HwMYPi7RSzXHO8wZaDdXgxN0u7tFxRV6H8OC1
ANTpOO6d6CFEIxuRIX6LXsQ3K0MTArU4IjNO7v5d/PTs6LT9dj+nMFA2njRBSOHaHUaZUqdPDlTZ
0jURIBf+Y2IyFMIyppMfOjkIwAl7OjnHetyt1iVz52r9Cy0f5G/3YWtWvxYXGP0eEIAWR3pTIsCC
ghrOtjgHzf4mI1BaVp5KK4l6MmSV0OZtC1IyGW6dyKcczcYPxXVDcIvKVG8BiXt422DppTKXommI
w3PSt+AtvAN1qb5SizokT9xhtzPpasm+imK3iaT0yGVvk/9VwZVGvpxetYBGt6aru9ahhNcrfIRz
tOs+O5ikxKeb9fva0l1AQKQnGyyzk/JRu/zbr8O2TmPFuwYuSfThCS32uoXE4O4O8T458UvYvI9o
AMaYjV3Hr99keCXWBOiHQL83XpUCXjIcVv3z9ZMVNm5FOIvJGPdYD08Ay174CIP7iabkjCD93/g4
Gs5N3DfmMOINbWDS5HiPBTqmQF8xL5P5uc0xp9wuoTXnNGxS4Hb2snPqb9wkg/Eui7f0YpDwbPPF
gG1mlHCO1iuPx1toJXVnM5VqGwaoCYYpAfj9QznmNTOHT7vA0q98Hp8GN3tEhbk3BsRiaWs8gu8X
BZpsRsHvC3aIh20RdZ9hyqagWp4Fnu71Rzfkbqn7weR8qn06ow4jKHR8XqUmihTODlX5rJ5wzP8F
sRbCbjborokfSoLTFjFpqKLIx17PERStmay18Ri2tBwyaK64t4FPJ95ZJ/aSqkaLoBpnC3R0E+cF
Ublq5AdTfotqhcoOA0onTMndP1AdMGGaUkYvbFb7+kBKfFwOkujtnGbYsT1xO5ay12z2vjm4h/mg
EI/bTXIS7l27AOjbz1PjUrw+jPttJLCryZI8loNOCIVwFiJ1gFsOjX1IiyeM5j295m0atFipURku
gT2sjBh1hfwpDH8NIqaqSYrSD1hJbCcNZpIUv2MoF+MtLaS4kA+BSP+4CQ9Af01bCRNnckbKUhUp
kjckiKlDSVnigGtoVTY333hR5wLk0YZlYLiNA2j/reyvhKzCEOUXMfFsTb3yUTyPrv2OhWsTug8w
/NhtL/QpVqfDUH9DKHcFa/XYwrnfsihV2odzP26ef2Gu/m+3aAH5TmQ30fx/mmJUjkSZQYoeQM/1
fFUhXVn2gpb0wPCq9YO21t4X7Y7TerH2o729ibyzfltqsipvUBAIIXNJ2kXs8k2sDQeoG4JQPp5O
ERGkqsufUy/E2n6UluXath7C3k3KzPkQELCeL+kJE+8zBUgRVQ1zdPkUfdAc6IHDSxT3vG6iO1YU
RXKkmjl7dT+DcPnh95b8hoeOcIF928U1tOFKhP0lwH4LDRF0VIb0QHTI9H/rXRBD+haxM+d32ril
lX34jAJrFi0D/vc/QCNlWNwSqYVT81aOPt/8FILZWOhiBey8en7xjILo3tSeIbqAcl3/SCFoNk89
qq8JOUP1dHgiqCXTnmivw3Xno8wdidaQpqgm1soJziD/tpgAnSKA62wxzUSAWcAofOB3PSRzgXq2
k0AynwjxPvfkDXuY8aDdYLWUHqnO0e1JdUoDdEoUrj0KScAujxrJNt0ZHGh0g597lXjLpRpZfJQ2
2pABbmKeLqbzXdRxH4W7pIQ13k6J1n+qxN2aTA98Vd7I4hL2GwYbf+1QObGqZAZhdzMTfXpTo2c4
r+h4/FMF+328BdSHGIsUNaXjblT6tpbxcVEtTEpMhawST5etqFGWbVHSeKG2npoRFBQ4VPtGnaDL
ha0LckJPVXOxjsDnZQXrbt+xw3BS7sugZfH6rInQjpTMB+0UBjArifL6W5SdZVq462RiMBoxrinH
4zEAl52+4Nqxz5BF/69Bsiht6pN1a398jyJsDy+cxlILh8MIBGJXP67QwzGMRjpacjQx5SwcrrJ3
Cj0pwlCyPNohLoM7XnCgKg8u/hxJeaUz/aKESa6AJTX3LZbXlFzJ7OQ9AoY1/SPPvaE1WwyMBfeK
C2U8GNhX1lOxBPvwc1vykulr/wjxbt6ZqGwYmrJyMspYBCHLtK8yPnAdIF8UgnPmH5qeW+dY62PP
utR4ezksKghPi0SCCUDus0JvFJ+pIJwna0uXCCCmzrG7epCUqkr3InuuX4lqypOEIowJcLBGnhwL
jFoF1Yhoz99W6NV0+PPZ3bgmiQzbD/iLlru7/PXsyZB8MhJUezUObJ1rBGKto2mIImGWdVZcr0FO
+L8msXUM9/AIog0ZlCSyD2Lf7jUfXYvg5HkCXcIYYh+orHnixYdz61owxRIn3USJBZI+0ckoKQ2w
yfaM8iUgdSGhCD57eXr25i9xM5yAqbFj+OJyStMCDb3iEO9jjkEJX0jGhUmHaKVeOLuYKyFsm/XO
rvsUBKmlXrmxVblvokBbcUpWWejp4g7sIU6fClJUc1oRE0V8coFCFJmod2KiTcsxNrY4RN4SRpC8
VDHOB2YEgnoFQkVndqTfgm/BrZ39gcWTXT8eQjGyQgd1grEwC6SqLsXqAj+tSPGpzWGs4xKpIJvS
SbiANbplKHhGMyugKGP1X/2VYKeUSyNEn7NWUDbpchTos9RVFZIFn1cb89PAx3K2OaIvPgA3lGln
1CYwKqG8GZudXArU2t1Et9iYcf37NJa/YqhzTi11JOs1xoib2Vu+Znw7a2d49laU3ZU7o8fXUuZ0
Q2w/a+Cf+VK1E84mE5j7+WJOkEW+xXAWuYZs6SfYDkd/w0kvfdyDm0a9/lp4endF4Hm3LIfyER/I
HrVDubfe1pBmEwzPIGmD3+M8y3d8vDeDe8Gm8cMDRijy8exifQNjkCehCxFlWtlavKXrVGYSWDx6
OohSxQzPjzN5X6J0ENpvwZQU5ocOqkktDHxlIWYCZndWZd3jXUskMTo36xEG/g9O3C0kpMVWAfKw
1dT7uqXlta0GpV2S9+W7A9TFGTZsbeeO1W1XJqwUg94sTF/DzUnvM+LkIA7YGiXSQczKQD5Q8lSI
GnFde5OK8Jxcw30vH/j/g2EFeJ9XH/vOgkxxFy8R9k/BPKq0mQWe5OG0YyupLU7xoYmJHSBUKiLO
9qQJxG/gS6LdWaYSNxPiMWF+C4W9un0+Uh7PT3hIAxtDRcwM3UCnjXyCODb4qxL2R4v/joWoKfcU
xB0zSwsvAJ1a+KYs3SwOKzMplUuHihm8J/GVnOfHKtL+J0JunTjLYDNLru77x2EYT8wyN7wCwDPN
MOss50cIwfrRT7GocudYBlutvXm24h4XM4+HG2pV8QmzJP4yzqv7WPf/TamuBsHn0XzszBspItSB
SE4+o6q7/cWg2QiZBg/sqHn9Oy3zryA4E5LXYYGIWKp9c845Ol/DqdsXgoHZvlAP+LC+vZ1ajOBH
PUivBI3O75E4Acjh35ymFke4AYnCbsdSO+IR/VK8keRkmQCDqbs4xfYcSPI0eeCUK9QfhsBHq2MD
N4pX066ofNTp1ktw4SFI3NDIToaSQfY09DHxAov07MhENR6Suk+dNJdatv7pMTXyVdpVhs09vj9b
Nw/HymZEfzzmNFvqeKbOfDQTvkKyK2iOSMktGAOKHeP78VxzmtR+GbDFoT8rV6yJCS/CJivIFLBz
OxcHVY+6tWTFHxPoSEAIrc+KNZnpC4lPNZX7kqfDDcpYtB+KkrnlnT+yziA9hhmMWw7OWwXw6+R7
jI1dgvp3GJ7aJmWc6xHVWNB5+a+ayofp3+vFb8FgpRIVPNIoQwV1pgCqJgM3uftVPgL8AsnAFY81
R4BeAUI17UhJAmmb1Yns+N7DR+cfS3XFCXOB8EtAfdr4JvFb+msnYVmSYhBebiV8kpkn0ZgWv+Ok
OtxdUmkavJ1kskqc057WjceraOdZ1vTMxfJeTZSIF6PaKKL4gSKjYenuqt/xztfHU7emPSbl3RRQ
qDqzZp5yYni9wMRzYTaT2fla86aKLxlCpqieEfiYtg1hSoJGq6mB0JugqS25E06CE67HKEw9Efp+
dplszzuAG48SZer4ghKfzfZOQ4BY4V3p/oeCcBUjCrlaQKeZA1xoQOWgbWvo9I8Imrlpp6fIUeZB
2a9Hb3pUGp/42tuvv48XAOXdDqmJ8ShEGzt/u+2jaY1VEwDeTgAhZqAaM/S6Gn9Ik67c2OMF2zLi
kKGtPMwPeSVcOKPMiCj+I+isTApNtpBQF+gy/wOd5MFhXMYsqcv0kigHIZ168FfRsS4dSslXmiY5
eYXyJpXBps0KIy6M9iZEmpXQXuw9BTr9Id0Vc6w7h9sfiBr7fZogW4DEnIBHmxIu692wo+aAWT9+
9Bb43cMOv1aRn6Qt1rR1qvLmoEmxsMKzS8LAjYsccalDKorsYelUDf/fv7BB7MNWQ6XIP7pI7uQF
6KxWHSH6bY1Cf3VFbTosYlUz0uOeLp3qAMuv1pY2fheW0gAdDBvCqlXrPTLCOksYxg1Ylfjv65jI
bly+OhuxtZreHrcUVr4cVAudvVFjFZYVnev+wipD7zOXZfPGPo//0lXZvMzez9mpywklyHf7c1Gw
W8KAyauBUCN3+U5G2TL6RdpnPtws9tJhMPlfbuRU8ZLiX+2rx/jdQsB4TjPVgHvRZ5cIlYlpRgvS
vMYu9IhJECR3yt+FqrFl7VR/RO8ph57UkBDvsccmaloB6XF2ZNMVy3V0+3YSduEpg3SE8ucCRO5M
LcANbH7oZ0GSrPaFYa0rZ6gXt6sUWaJ4UUAQDBI69rZEOBBEJUKEmXgtkuzgsGplAGS0aP8DPjMc
WHdMTNtQIwA3qz0pc+eyU9KMMcOihmRVo6v05CfMMchb/2rDcx702l+qIt07Dx5igWDJo8Ba62/5
G88h0s/b2x6XyUA/3BMuMI8vkzYxrrAq2XtwLx7LBlnKTSZs7JoAQ+7nS6XeGYf747T2ZONSB1qW
ZgA7CeDNM+39WsKfwGnnuXYrGSh3YnWTgurKScDKM0PBk5uj6yBiyNXjPF9S8i1c7rXscVpiZ0gU
c4lT/LcUNaQ96aBK0x4IY6eZNew+85f4mcjzV/w/no99oabvNedOkilb6lz3t5KtLfp3cU3XUST2
k0yFhLeTHkKc014FAgkfd7N+KNBaVH156mUGcmY9hPIg8UKwoGXPpiFuDa2/Sj2uqCmvixvYvlkg
s8DVzYUQlHydSU4HKe5r47612Dc1QQd2Dn/w6KCTJ5+AF/0Ru2/EASTZ8oiZSiUoFQT5Nzt5Zbmf
PqzJHbOJQFL3HtO01AuFFwVX+ff0YAy63380CJVIGguZWlM//+dAiQJnnc7P7nApIG30Fx55sA3y
KyxA9cwfM52QpS4w5zOKQHlKzt3d+nVGFHggzO9bXYKgqWvW/qay+44B5XP+vDHt0NirnYX4nasE
ptiGHPQ3EQWnWcBS8Mlhi/fuAqv2UPEXXP5UmC3u0WRfTaPhJOdLqtJCG0hlcfc6oR7A7bYP0ciz
+tm2jKCcTaIahmUUNvzZAUUZjhXtKG5q5ven+RYq1MG4rjx++FBSQaZ2+aOPqYbuK5efoQOCwmuD
Osj5KfeXckPw3Ocv0crf9C//PnxCRJz2L5hqZ7G2v9aS4+rVAt95/f1P2VH0vkVZ6TqRDsxK1+4l
3BlAn8tq3MXaQYs1
`protect end_protected
